// Generator : SpinalHDL v1.9.4    git head : 270018552577f3bb8e5339ee2583c9c22d324215
// Component : NV_NVDLA_CDMA_shared_buffer
// Git hash  : e8247006974f01f499a02b4ce7fad5c2ba9dc983

`timescale 1ns/1ps

module NV_NVDLA_CDMA_shared_buffer (
  input  wire          dc2sbuf_p_wr_0_addr_valid,
  input  wire [7:0]    dc2sbuf_p_wr_0_addr_payload,
  input  wire [63:0]   dc2sbuf_p_wr_0_data,
  input  wire          dc2sbuf_p_wr_1_addr_valid,
  input  wire [7:0]    dc2sbuf_p_wr_1_addr_payload,
  input  wire [63:0]   dc2sbuf_p_wr_1_data,
  input  wire          img2sbuf_p_wr_0_addr_valid,
  input  wire [7:0]    img2sbuf_p_wr_0_addr_payload,
  input  wire [63:0]   img2sbuf_p_wr_0_data,
  input  wire          img2sbuf_p_wr_1_addr_valid,
  input  wire [7:0]    img2sbuf_p_wr_1_addr_payload,
  input  wire [63:0]   img2sbuf_p_wr_1_data,
  input  wire          dc2sbuf_p_rd_0_addr_valid,
  input  wire [7:0]    dc2sbuf_p_rd_0_addr_payload,
  output wire [63:0]   dc2sbuf_p_rd_0_data,
  input  wire          dc2sbuf_p_rd_1_addr_valid,
  input  wire [7:0]    dc2sbuf_p_rd_1_addr_payload,
  output wire [63:0]   dc2sbuf_p_rd_1_data,
  input  wire          img2sbuf_p_rd_0_addr_valid,
  input  wire [7:0]    img2sbuf_p_rd_0_addr_payload,
  output wire [63:0]   img2sbuf_p_rd_0_data,
  input  wire          img2sbuf_p_rd_1_addr_valid,
  input  wire [7:0]    img2sbuf_p_rd_1_addr_payload,
  output wire [63:0]   img2sbuf_p_rd_1_data,
  input  wire          clk,
  input  wire          reset
);

  wire       [63:0]   shareBuffer_buffer_0_dout;
  wire       [63:0]   shareBuffer_buffer_1_dout;
  wire       [63:0]   shareBuffer_buffer_2_dout;
  wire       [63:0]   shareBuffer_buffer_3_dout;
  wire       [63:0]   shareBuffer_buffer_4_dout;
  wire       [63:0]   shareBuffer_buffer_5_dout;
  wire       [63:0]   shareBuffer_buffer_6_dout;
  wire       [63:0]   shareBuffer_buffer_7_dout;
  wire       [63:0]   shareBuffer_buffer_8_dout;
  wire       [63:0]   shareBuffer_buffer_9_dout;
  wire       [63:0]   shareBuffer_buffer_10_dout;
  wire       [63:0]   shareBuffer_buffer_11_dout;
  wire       [63:0]   shareBuffer_buffer_12_dout;
  wire       [63:0]   shareBuffer_buffer_13_dout;
  wire       [63:0]   shareBuffer_buffer_14_dout;
  wire       [63:0]   shareBuffer_buffer_15_dout;
  wire       [0:0]    _zz_sbuf_wa_0;
  wire       [2:0]    _zz_sbuf_wa_0_1;
  wire       [3:0]    _zz_sbuf_wa_0_2;
  wire       [0:0]    _zz_sbuf_wa_0_3;
  wire       [2:0]    _zz_sbuf_wa_0_4;
  wire       [3:0]    _zz_sbuf_wa_0_5;
  wire       [0:0]    _zz_sbuf_wa_0_6;
  wire       [1:0]    _zz_sbuf_wa_0_7;
  wire       [0:0]    _zz_sbuf_wa_0_8;
  wire       [0:0]    _zz_sbuf_wa_0_9;
  wire       [0:0]    _zz_sbuf_wa_1;
  wire       [2:0]    _zz_sbuf_wa_1_1;
  wire       [3:0]    _zz_sbuf_wa_1_2;
  wire       [0:0]    _zz_sbuf_wa_1_3;
  wire       [2:0]    _zz_sbuf_wa_1_4;
  wire       [3:0]    _zz_sbuf_wa_1_5;
  wire       [0:0]    _zz_sbuf_wa_1_6;
  wire       [1:0]    _zz_sbuf_wa_1_7;
  wire       [0:0]    _zz_sbuf_wa_1_8;
  wire       [0:0]    _zz_sbuf_wa_1_9;
  wire       [0:0]    _zz_sbuf_wa_2;
  wire       [2:0]    _zz_sbuf_wa_2_1;
  wire       [3:0]    _zz_sbuf_wa_2_2;
  wire       [0:0]    _zz_sbuf_wa_2_3;
  wire       [2:0]    _zz_sbuf_wa_2_4;
  wire       [3:0]    _zz_sbuf_wa_2_5;
  wire       [0:0]    _zz_sbuf_wa_2_6;
  wire       [1:0]    _zz_sbuf_wa_2_7;
  wire       [0:0]    _zz_sbuf_wa_2_8;
  wire       [0:0]    _zz_sbuf_wa_2_9;
  wire       [0:0]    _zz_sbuf_wa_3;
  wire       [2:0]    _zz_sbuf_wa_3_1;
  wire       [3:0]    _zz_sbuf_wa_3_2;
  wire       [0:0]    _zz_sbuf_wa_3_3;
  wire       [2:0]    _zz_sbuf_wa_3_4;
  wire       [3:0]    _zz_sbuf_wa_3_5;
  wire       [0:0]    _zz_sbuf_wa_3_6;
  wire       [1:0]    _zz_sbuf_wa_3_7;
  wire       [0:0]    _zz_sbuf_wa_3_8;
  wire       [0:0]    _zz_sbuf_wa_3_9;
  wire       [0:0]    _zz_sbuf_wa_4;
  wire       [2:0]    _zz_sbuf_wa_4_1;
  wire       [3:0]    _zz_sbuf_wa_4_2;
  wire       [0:0]    _zz_sbuf_wa_4_3;
  wire       [2:0]    _zz_sbuf_wa_4_4;
  wire       [3:0]    _zz_sbuf_wa_4_5;
  wire       [0:0]    _zz_sbuf_wa_4_6;
  wire       [1:0]    _zz_sbuf_wa_4_7;
  wire       [0:0]    _zz_sbuf_wa_4_8;
  wire       [0:0]    _zz_sbuf_wa_4_9;
  wire       [0:0]    _zz_sbuf_wa_5;
  wire       [2:0]    _zz_sbuf_wa_5_1;
  wire       [3:0]    _zz_sbuf_wa_5_2;
  wire       [0:0]    _zz_sbuf_wa_5_3;
  wire       [2:0]    _zz_sbuf_wa_5_4;
  wire       [3:0]    _zz_sbuf_wa_5_5;
  wire       [0:0]    _zz_sbuf_wa_5_6;
  wire       [1:0]    _zz_sbuf_wa_5_7;
  wire       [0:0]    _zz_sbuf_wa_5_8;
  wire       [0:0]    _zz_sbuf_wa_5_9;
  wire       [0:0]    _zz_sbuf_wa_6;
  wire       [2:0]    _zz_sbuf_wa_6_1;
  wire       [3:0]    _zz_sbuf_wa_6_2;
  wire       [0:0]    _zz_sbuf_wa_6_3;
  wire       [2:0]    _zz_sbuf_wa_6_4;
  wire       [3:0]    _zz_sbuf_wa_6_5;
  wire       [0:0]    _zz_sbuf_wa_6_6;
  wire       [1:0]    _zz_sbuf_wa_6_7;
  wire       [0:0]    _zz_sbuf_wa_6_8;
  wire       [0:0]    _zz_sbuf_wa_6_9;
  wire       [0:0]    _zz_sbuf_wa_7;
  wire       [2:0]    _zz_sbuf_wa_7_1;
  wire       [3:0]    _zz_sbuf_wa_7_2;
  wire       [0:0]    _zz_sbuf_wa_7_3;
  wire       [2:0]    _zz_sbuf_wa_7_4;
  wire       [3:0]    _zz_sbuf_wa_7_5;
  wire       [0:0]    _zz_sbuf_wa_7_6;
  wire       [1:0]    _zz_sbuf_wa_7_7;
  wire       [0:0]    _zz_sbuf_wa_7_8;
  wire       [0:0]    _zz_sbuf_wa_7_9;
  wire       [0:0]    _zz_sbuf_wa_8;
  wire       [2:0]    _zz_sbuf_wa_8_1;
  wire       [3:0]    _zz_sbuf_wa_8_2;
  wire       [0:0]    _zz_sbuf_wa_8_3;
  wire       [2:0]    _zz_sbuf_wa_8_4;
  wire       [3:0]    _zz_sbuf_wa_8_5;
  wire       [0:0]    _zz_sbuf_wa_8_6;
  wire       [1:0]    _zz_sbuf_wa_8_7;
  wire       [0:0]    _zz_sbuf_wa_8_8;
  wire       [0:0]    _zz_sbuf_wa_8_9;
  wire       [0:0]    _zz_sbuf_wa_9;
  wire       [2:0]    _zz_sbuf_wa_9_1;
  wire       [3:0]    _zz_sbuf_wa_9_2;
  wire       [0:0]    _zz_sbuf_wa_9_3;
  wire       [2:0]    _zz_sbuf_wa_9_4;
  wire       [3:0]    _zz_sbuf_wa_9_5;
  wire       [0:0]    _zz_sbuf_wa_9_6;
  wire       [1:0]    _zz_sbuf_wa_9_7;
  wire       [0:0]    _zz_sbuf_wa_9_8;
  wire       [0:0]    _zz_sbuf_wa_9_9;
  wire       [0:0]    _zz_sbuf_wa_10;
  wire       [2:0]    _zz_sbuf_wa_10_1;
  wire       [3:0]    _zz_sbuf_wa_10_2;
  wire       [0:0]    _zz_sbuf_wa_10_3;
  wire       [2:0]    _zz_sbuf_wa_10_4;
  wire       [3:0]    _zz_sbuf_wa_10_5;
  wire       [0:0]    _zz_sbuf_wa_10_6;
  wire       [1:0]    _zz_sbuf_wa_10_7;
  wire       [0:0]    _zz_sbuf_wa_10_8;
  wire       [0:0]    _zz_sbuf_wa_10_9;
  wire       [0:0]    _zz_sbuf_wa_11;
  wire       [2:0]    _zz_sbuf_wa_11_1;
  wire       [3:0]    _zz_sbuf_wa_11_2;
  wire       [0:0]    _zz_sbuf_wa_11_3;
  wire       [2:0]    _zz_sbuf_wa_11_4;
  wire       [3:0]    _zz_sbuf_wa_11_5;
  wire       [0:0]    _zz_sbuf_wa_11_6;
  wire       [1:0]    _zz_sbuf_wa_11_7;
  wire       [0:0]    _zz_sbuf_wa_11_8;
  wire       [0:0]    _zz_sbuf_wa_11_9;
  wire       [0:0]    _zz_sbuf_wa_12;
  wire       [2:0]    _zz_sbuf_wa_12_1;
  wire       [3:0]    _zz_sbuf_wa_12_2;
  wire       [0:0]    _zz_sbuf_wa_12_3;
  wire       [2:0]    _zz_sbuf_wa_12_4;
  wire       [3:0]    _zz_sbuf_wa_12_5;
  wire       [0:0]    _zz_sbuf_wa_12_6;
  wire       [1:0]    _zz_sbuf_wa_12_7;
  wire       [0:0]    _zz_sbuf_wa_12_8;
  wire       [0:0]    _zz_sbuf_wa_12_9;
  wire       [0:0]    _zz_sbuf_wa_13;
  wire       [2:0]    _zz_sbuf_wa_13_1;
  wire       [3:0]    _zz_sbuf_wa_13_2;
  wire       [0:0]    _zz_sbuf_wa_13_3;
  wire       [2:0]    _zz_sbuf_wa_13_4;
  wire       [3:0]    _zz_sbuf_wa_13_5;
  wire       [0:0]    _zz_sbuf_wa_13_6;
  wire       [1:0]    _zz_sbuf_wa_13_7;
  wire       [0:0]    _zz_sbuf_wa_13_8;
  wire       [0:0]    _zz_sbuf_wa_13_9;
  wire       [0:0]    _zz_sbuf_wa_14;
  wire       [2:0]    _zz_sbuf_wa_14_1;
  wire       [3:0]    _zz_sbuf_wa_14_2;
  wire       [0:0]    _zz_sbuf_wa_14_3;
  wire       [2:0]    _zz_sbuf_wa_14_4;
  wire       [3:0]    _zz_sbuf_wa_14_5;
  wire       [0:0]    _zz_sbuf_wa_14_6;
  wire       [1:0]    _zz_sbuf_wa_14_7;
  wire       [0:0]    _zz_sbuf_wa_14_8;
  wire       [0:0]    _zz_sbuf_wa_14_9;
  wire       [0:0]    _zz_sbuf_wa_15;
  wire       [2:0]    _zz_sbuf_wa_15_1;
  wire       [3:0]    _zz_sbuf_wa_15_2;
  wire       [0:0]    _zz_sbuf_wa_15_3;
  wire       [2:0]    _zz_sbuf_wa_15_4;
  wire       [3:0]    _zz_sbuf_wa_15_5;
  wire       [0:0]    _zz_sbuf_wa_15_6;
  wire       [1:0]    _zz_sbuf_wa_15_7;
  wire       [0:0]    _zz_sbuf_wa_15_8;
  wire       [0:0]    _zz_sbuf_wa_15_9;
  wire       [0:0]    _zz_sbuf_wdat_0;
  wire       [61:0]   _zz_sbuf_wdat_0_1;
  wire       [0:0]    _zz_sbuf_wdat_0_2;
  wire       [57:0]   _zz_sbuf_wdat_0_3;
  wire       [0:0]    _zz_sbuf_wdat_0_4;
  wire       [53:0]   _zz_sbuf_wdat_0_5;
  wire       [0:0]    _zz_sbuf_wdat_0_6;
  wire       [49:0]   _zz_sbuf_wdat_0_7;
  wire       [0:0]    _zz_sbuf_wdat_0_8;
  wire       [45:0]   _zz_sbuf_wdat_0_9;
  wire       [0:0]    _zz_sbuf_wdat_0_10;
  wire       [41:0]   _zz_sbuf_wdat_0_11;
  wire       [0:0]    _zz_sbuf_wdat_0_12;
  wire       [37:0]   _zz_sbuf_wdat_0_13;
  wire       [0:0]    _zz_sbuf_wdat_0_14;
  wire       [33:0]   _zz_sbuf_wdat_0_15;
  wire       [0:0]    _zz_sbuf_wdat_0_16;
  wire       [29:0]   _zz_sbuf_wdat_0_17;
  wire       [0:0]    _zz_sbuf_wdat_0_18;
  wire       [25:0]   _zz_sbuf_wdat_0_19;
  wire       [0:0]    _zz_sbuf_wdat_0_20;
  wire       [21:0]   _zz_sbuf_wdat_0_21;
  wire       [0:0]    _zz_sbuf_wdat_0_22;
  wire       [17:0]   _zz_sbuf_wdat_0_23;
  wire       [0:0]    _zz_sbuf_wdat_0_24;
  wire       [13:0]   _zz_sbuf_wdat_0_25;
  wire       [0:0]    _zz_sbuf_wdat_0_26;
  wire       [9:0]    _zz_sbuf_wdat_0_27;
  wire       [0:0]    _zz_sbuf_wdat_0_28;
  wire       [5:0]    _zz_sbuf_wdat_0_29;
  wire       [0:0]    _zz_sbuf_wdat_0_30;
  wire       [0:0]    _zz_sbuf_wdat_0_31;
  wire       [0:0]    _zz_sbuf_wdat_0_32;
  wire       [61:0]   _zz_sbuf_wdat_0_33;
  wire       [0:0]    _zz_sbuf_wdat_0_34;
  wire       [57:0]   _zz_sbuf_wdat_0_35;
  wire       [0:0]    _zz_sbuf_wdat_0_36;
  wire       [53:0]   _zz_sbuf_wdat_0_37;
  wire       [0:0]    _zz_sbuf_wdat_0_38;
  wire       [49:0]   _zz_sbuf_wdat_0_39;
  wire       [0:0]    _zz_sbuf_wdat_0_40;
  wire       [45:0]   _zz_sbuf_wdat_0_41;
  wire       [0:0]    _zz_sbuf_wdat_0_42;
  wire       [41:0]   _zz_sbuf_wdat_0_43;
  wire       [0:0]    _zz_sbuf_wdat_0_44;
  wire       [37:0]   _zz_sbuf_wdat_0_45;
  wire       [0:0]    _zz_sbuf_wdat_0_46;
  wire       [33:0]   _zz_sbuf_wdat_0_47;
  wire       [0:0]    _zz_sbuf_wdat_0_48;
  wire       [29:0]   _zz_sbuf_wdat_0_49;
  wire       [0:0]    _zz_sbuf_wdat_0_50;
  wire       [25:0]   _zz_sbuf_wdat_0_51;
  wire       [0:0]    _zz_sbuf_wdat_0_52;
  wire       [21:0]   _zz_sbuf_wdat_0_53;
  wire       [0:0]    _zz_sbuf_wdat_0_54;
  wire       [17:0]   _zz_sbuf_wdat_0_55;
  wire       [0:0]    _zz_sbuf_wdat_0_56;
  wire       [13:0]   _zz_sbuf_wdat_0_57;
  wire       [0:0]    _zz_sbuf_wdat_0_58;
  wire       [9:0]    _zz_sbuf_wdat_0_59;
  wire       [0:0]    _zz_sbuf_wdat_0_60;
  wire       [5:0]    _zz_sbuf_wdat_0_61;
  wire       [0:0]    _zz_sbuf_wdat_0_62;
  wire       [0:0]    _zz_sbuf_wdat_0_63;
  wire       [0:0]    _zz_sbuf_wdat_0_64;
  wire       [60:0]   _zz_sbuf_wdat_0_65;
  wire       [0:0]    _zz_sbuf_wdat_0_66;
  wire       [56:0]   _zz_sbuf_wdat_0_67;
  wire       [0:0]    _zz_sbuf_wdat_0_68;
  wire       [52:0]   _zz_sbuf_wdat_0_69;
  wire       [0:0]    _zz_sbuf_wdat_0_70;
  wire       [48:0]   _zz_sbuf_wdat_0_71;
  wire       [0:0]    _zz_sbuf_wdat_0_72;
  wire       [44:0]   _zz_sbuf_wdat_0_73;
  wire       [0:0]    _zz_sbuf_wdat_0_74;
  wire       [40:0]   _zz_sbuf_wdat_0_75;
  wire       [0:0]    _zz_sbuf_wdat_0_76;
  wire       [36:0]   _zz_sbuf_wdat_0_77;
  wire       [0:0]    _zz_sbuf_wdat_0_78;
  wire       [32:0]   _zz_sbuf_wdat_0_79;
  wire       [0:0]    _zz_sbuf_wdat_0_80;
  wire       [28:0]   _zz_sbuf_wdat_0_81;
  wire       [0:0]    _zz_sbuf_wdat_0_82;
  wire       [24:0]   _zz_sbuf_wdat_0_83;
  wire       [0:0]    _zz_sbuf_wdat_0_84;
  wire       [20:0]   _zz_sbuf_wdat_0_85;
  wire       [0:0]    _zz_sbuf_wdat_0_86;
  wire       [16:0]   _zz_sbuf_wdat_0_87;
  wire       [0:0]    _zz_sbuf_wdat_0_88;
  wire       [12:0]   _zz_sbuf_wdat_0_89;
  wire       [0:0]    _zz_sbuf_wdat_0_90;
  wire       [8:0]    _zz_sbuf_wdat_0_91;
  wire       [0:0]    _zz_sbuf_wdat_0_92;
  wire       [4:0]    _zz_sbuf_wdat_0_93;
  wire       [0:0]    _zz_sbuf_wdat_0_94;
  wire       [59:0]   _zz_sbuf_wdat_0_95;
  wire       [0:0]    _zz_sbuf_wdat_0_96;
  wire       [55:0]   _zz_sbuf_wdat_0_97;
  wire       [0:0]    _zz_sbuf_wdat_0_98;
  wire       [51:0]   _zz_sbuf_wdat_0_99;
  wire       [0:0]    _zz_sbuf_wdat_0_100;
  wire       [47:0]   _zz_sbuf_wdat_0_101;
  wire       [0:0]    _zz_sbuf_wdat_0_102;
  wire       [43:0]   _zz_sbuf_wdat_0_103;
  wire       [0:0]    _zz_sbuf_wdat_0_104;
  wire       [39:0]   _zz_sbuf_wdat_0_105;
  wire       [0:0]    _zz_sbuf_wdat_0_106;
  wire       [35:0]   _zz_sbuf_wdat_0_107;
  wire       [0:0]    _zz_sbuf_wdat_0_108;
  wire       [31:0]   _zz_sbuf_wdat_0_109;
  wire       [0:0]    _zz_sbuf_wdat_0_110;
  wire       [27:0]   _zz_sbuf_wdat_0_111;
  wire       [0:0]    _zz_sbuf_wdat_0_112;
  wire       [23:0]   _zz_sbuf_wdat_0_113;
  wire       [0:0]    _zz_sbuf_wdat_0_114;
  wire       [19:0]   _zz_sbuf_wdat_0_115;
  wire       [0:0]    _zz_sbuf_wdat_0_116;
  wire       [15:0]   _zz_sbuf_wdat_0_117;
  wire       [0:0]    _zz_sbuf_wdat_0_118;
  wire       [11:0]   _zz_sbuf_wdat_0_119;
  wire       [0:0]    _zz_sbuf_wdat_0_120;
  wire       [7:0]    _zz_sbuf_wdat_0_121;
  wire       [0:0]    _zz_sbuf_wdat_0_122;
  wire       [3:0]    _zz_sbuf_wdat_0_123;
  wire       [0:0]    _zz_sbuf_wdat_1;
  wire       [61:0]   _zz_sbuf_wdat_1_1;
  wire       [0:0]    _zz_sbuf_wdat_1_2;
  wire       [57:0]   _zz_sbuf_wdat_1_3;
  wire       [0:0]    _zz_sbuf_wdat_1_4;
  wire       [53:0]   _zz_sbuf_wdat_1_5;
  wire       [0:0]    _zz_sbuf_wdat_1_6;
  wire       [49:0]   _zz_sbuf_wdat_1_7;
  wire       [0:0]    _zz_sbuf_wdat_1_8;
  wire       [45:0]   _zz_sbuf_wdat_1_9;
  wire       [0:0]    _zz_sbuf_wdat_1_10;
  wire       [41:0]   _zz_sbuf_wdat_1_11;
  wire       [0:0]    _zz_sbuf_wdat_1_12;
  wire       [37:0]   _zz_sbuf_wdat_1_13;
  wire       [0:0]    _zz_sbuf_wdat_1_14;
  wire       [33:0]   _zz_sbuf_wdat_1_15;
  wire       [0:0]    _zz_sbuf_wdat_1_16;
  wire       [29:0]   _zz_sbuf_wdat_1_17;
  wire       [0:0]    _zz_sbuf_wdat_1_18;
  wire       [25:0]   _zz_sbuf_wdat_1_19;
  wire       [0:0]    _zz_sbuf_wdat_1_20;
  wire       [21:0]   _zz_sbuf_wdat_1_21;
  wire       [0:0]    _zz_sbuf_wdat_1_22;
  wire       [17:0]   _zz_sbuf_wdat_1_23;
  wire       [0:0]    _zz_sbuf_wdat_1_24;
  wire       [13:0]   _zz_sbuf_wdat_1_25;
  wire       [0:0]    _zz_sbuf_wdat_1_26;
  wire       [9:0]    _zz_sbuf_wdat_1_27;
  wire       [0:0]    _zz_sbuf_wdat_1_28;
  wire       [5:0]    _zz_sbuf_wdat_1_29;
  wire       [0:0]    _zz_sbuf_wdat_1_30;
  wire       [0:0]    _zz_sbuf_wdat_1_31;
  wire       [0:0]    _zz_sbuf_wdat_1_32;
  wire       [61:0]   _zz_sbuf_wdat_1_33;
  wire       [0:0]    _zz_sbuf_wdat_1_34;
  wire       [57:0]   _zz_sbuf_wdat_1_35;
  wire       [0:0]    _zz_sbuf_wdat_1_36;
  wire       [53:0]   _zz_sbuf_wdat_1_37;
  wire       [0:0]    _zz_sbuf_wdat_1_38;
  wire       [49:0]   _zz_sbuf_wdat_1_39;
  wire       [0:0]    _zz_sbuf_wdat_1_40;
  wire       [45:0]   _zz_sbuf_wdat_1_41;
  wire       [0:0]    _zz_sbuf_wdat_1_42;
  wire       [41:0]   _zz_sbuf_wdat_1_43;
  wire       [0:0]    _zz_sbuf_wdat_1_44;
  wire       [37:0]   _zz_sbuf_wdat_1_45;
  wire       [0:0]    _zz_sbuf_wdat_1_46;
  wire       [33:0]   _zz_sbuf_wdat_1_47;
  wire       [0:0]    _zz_sbuf_wdat_1_48;
  wire       [29:0]   _zz_sbuf_wdat_1_49;
  wire       [0:0]    _zz_sbuf_wdat_1_50;
  wire       [25:0]   _zz_sbuf_wdat_1_51;
  wire       [0:0]    _zz_sbuf_wdat_1_52;
  wire       [21:0]   _zz_sbuf_wdat_1_53;
  wire       [0:0]    _zz_sbuf_wdat_1_54;
  wire       [17:0]   _zz_sbuf_wdat_1_55;
  wire       [0:0]    _zz_sbuf_wdat_1_56;
  wire       [13:0]   _zz_sbuf_wdat_1_57;
  wire       [0:0]    _zz_sbuf_wdat_1_58;
  wire       [9:0]    _zz_sbuf_wdat_1_59;
  wire       [0:0]    _zz_sbuf_wdat_1_60;
  wire       [5:0]    _zz_sbuf_wdat_1_61;
  wire       [0:0]    _zz_sbuf_wdat_1_62;
  wire       [0:0]    _zz_sbuf_wdat_1_63;
  wire       [0:0]    _zz_sbuf_wdat_1_64;
  wire       [60:0]   _zz_sbuf_wdat_1_65;
  wire       [0:0]    _zz_sbuf_wdat_1_66;
  wire       [56:0]   _zz_sbuf_wdat_1_67;
  wire       [0:0]    _zz_sbuf_wdat_1_68;
  wire       [52:0]   _zz_sbuf_wdat_1_69;
  wire       [0:0]    _zz_sbuf_wdat_1_70;
  wire       [48:0]   _zz_sbuf_wdat_1_71;
  wire       [0:0]    _zz_sbuf_wdat_1_72;
  wire       [44:0]   _zz_sbuf_wdat_1_73;
  wire       [0:0]    _zz_sbuf_wdat_1_74;
  wire       [40:0]   _zz_sbuf_wdat_1_75;
  wire       [0:0]    _zz_sbuf_wdat_1_76;
  wire       [36:0]   _zz_sbuf_wdat_1_77;
  wire       [0:0]    _zz_sbuf_wdat_1_78;
  wire       [32:0]   _zz_sbuf_wdat_1_79;
  wire       [0:0]    _zz_sbuf_wdat_1_80;
  wire       [28:0]   _zz_sbuf_wdat_1_81;
  wire       [0:0]    _zz_sbuf_wdat_1_82;
  wire       [24:0]   _zz_sbuf_wdat_1_83;
  wire       [0:0]    _zz_sbuf_wdat_1_84;
  wire       [20:0]   _zz_sbuf_wdat_1_85;
  wire       [0:0]    _zz_sbuf_wdat_1_86;
  wire       [16:0]   _zz_sbuf_wdat_1_87;
  wire       [0:0]    _zz_sbuf_wdat_1_88;
  wire       [12:0]   _zz_sbuf_wdat_1_89;
  wire       [0:0]    _zz_sbuf_wdat_1_90;
  wire       [8:0]    _zz_sbuf_wdat_1_91;
  wire       [0:0]    _zz_sbuf_wdat_1_92;
  wire       [4:0]    _zz_sbuf_wdat_1_93;
  wire       [0:0]    _zz_sbuf_wdat_1_94;
  wire       [59:0]   _zz_sbuf_wdat_1_95;
  wire       [0:0]    _zz_sbuf_wdat_1_96;
  wire       [55:0]   _zz_sbuf_wdat_1_97;
  wire       [0:0]    _zz_sbuf_wdat_1_98;
  wire       [51:0]   _zz_sbuf_wdat_1_99;
  wire       [0:0]    _zz_sbuf_wdat_1_100;
  wire       [47:0]   _zz_sbuf_wdat_1_101;
  wire       [0:0]    _zz_sbuf_wdat_1_102;
  wire       [43:0]   _zz_sbuf_wdat_1_103;
  wire       [0:0]    _zz_sbuf_wdat_1_104;
  wire       [39:0]   _zz_sbuf_wdat_1_105;
  wire       [0:0]    _zz_sbuf_wdat_1_106;
  wire       [35:0]   _zz_sbuf_wdat_1_107;
  wire       [0:0]    _zz_sbuf_wdat_1_108;
  wire       [31:0]   _zz_sbuf_wdat_1_109;
  wire       [0:0]    _zz_sbuf_wdat_1_110;
  wire       [27:0]   _zz_sbuf_wdat_1_111;
  wire       [0:0]    _zz_sbuf_wdat_1_112;
  wire       [23:0]   _zz_sbuf_wdat_1_113;
  wire       [0:0]    _zz_sbuf_wdat_1_114;
  wire       [19:0]   _zz_sbuf_wdat_1_115;
  wire       [0:0]    _zz_sbuf_wdat_1_116;
  wire       [15:0]   _zz_sbuf_wdat_1_117;
  wire       [0:0]    _zz_sbuf_wdat_1_118;
  wire       [11:0]   _zz_sbuf_wdat_1_119;
  wire       [0:0]    _zz_sbuf_wdat_1_120;
  wire       [7:0]    _zz_sbuf_wdat_1_121;
  wire       [0:0]    _zz_sbuf_wdat_1_122;
  wire       [3:0]    _zz_sbuf_wdat_1_123;
  wire       [0:0]    _zz_sbuf_wdat_2;
  wire       [61:0]   _zz_sbuf_wdat_2_1;
  wire       [0:0]    _zz_sbuf_wdat_2_2;
  wire       [57:0]   _zz_sbuf_wdat_2_3;
  wire       [0:0]    _zz_sbuf_wdat_2_4;
  wire       [53:0]   _zz_sbuf_wdat_2_5;
  wire       [0:0]    _zz_sbuf_wdat_2_6;
  wire       [49:0]   _zz_sbuf_wdat_2_7;
  wire       [0:0]    _zz_sbuf_wdat_2_8;
  wire       [45:0]   _zz_sbuf_wdat_2_9;
  wire       [0:0]    _zz_sbuf_wdat_2_10;
  wire       [41:0]   _zz_sbuf_wdat_2_11;
  wire       [0:0]    _zz_sbuf_wdat_2_12;
  wire       [37:0]   _zz_sbuf_wdat_2_13;
  wire       [0:0]    _zz_sbuf_wdat_2_14;
  wire       [33:0]   _zz_sbuf_wdat_2_15;
  wire       [0:0]    _zz_sbuf_wdat_2_16;
  wire       [29:0]   _zz_sbuf_wdat_2_17;
  wire       [0:0]    _zz_sbuf_wdat_2_18;
  wire       [25:0]   _zz_sbuf_wdat_2_19;
  wire       [0:0]    _zz_sbuf_wdat_2_20;
  wire       [21:0]   _zz_sbuf_wdat_2_21;
  wire       [0:0]    _zz_sbuf_wdat_2_22;
  wire       [17:0]   _zz_sbuf_wdat_2_23;
  wire       [0:0]    _zz_sbuf_wdat_2_24;
  wire       [13:0]   _zz_sbuf_wdat_2_25;
  wire       [0:0]    _zz_sbuf_wdat_2_26;
  wire       [9:0]    _zz_sbuf_wdat_2_27;
  wire       [0:0]    _zz_sbuf_wdat_2_28;
  wire       [5:0]    _zz_sbuf_wdat_2_29;
  wire       [0:0]    _zz_sbuf_wdat_2_30;
  wire       [0:0]    _zz_sbuf_wdat_2_31;
  wire       [0:0]    _zz_sbuf_wdat_2_32;
  wire       [61:0]   _zz_sbuf_wdat_2_33;
  wire       [0:0]    _zz_sbuf_wdat_2_34;
  wire       [57:0]   _zz_sbuf_wdat_2_35;
  wire       [0:0]    _zz_sbuf_wdat_2_36;
  wire       [53:0]   _zz_sbuf_wdat_2_37;
  wire       [0:0]    _zz_sbuf_wdat_2_38;
  wire       [49:0]   _zz_sbuf_wdat_2_39;
  wire       [0:0]    _zz_sbuf_wdat_2_40;
  wire       [45:0]   _zz_sbuf_wdat_2_41;
  wire       [0:0]    _zz_sbuf_wdat_2_42;
  wire       [41:0]   _zz_sbuf_wdat_2_43;
  wire       [0:0]    _zz_sbuf_wdat_2_44;
  wire       [37:0]   _zz_sbuf_wdat_2_45;
  wire       [0:0]    _zz_sbuf_wdat_2_46;
  wire       [33:0]   _zz_sbuf_wdat_2_47;
  wire       [0:0]    _zz_sbuf_wdat_2_48;
  wire       [29:0]   _zz_sbuf_wdat_2_49;
  wire       [0:0]    _zz_sbuf_wdat_2_50;
  wire       [25:0]   _zz_sbuf_wdat_2_51;
  wire       [0:0]    _zz_sbuf_wdat_2_52;
  wire       [21:0]   _zz_sbuf_wdat_2_53;
  wire       [0:0]    _zz_sbuf_wdat_2_54;
  wire       [17:0]   _zz_sbuf_wdat_2_55;
  wire       [0:0]    _zz_sbuf_wdat_2_56;
  wire       [13:0]   _zz_sbuf_wdat_2_57;
  wire       [0:0]    _zz_sbuf_wdat_2_58;
  wire       [9:0]    _zz_sbuf_wdat_2_59;
  wire       [0:0]    _zz_sbuf_wdat_2_60;
  wire       [5:0]    _zz_sbuf_wdat_2_61;
  wire       [0:0]    _zz_sbuf_wdat_2_62;
  wire       [0:0]    _zz_sbuf_wdat_2_63;
  wire       [0:0]    _zz_sbuf_wdat_2_64;
  wire       [60:0]   _zz_sbuf_wdat_2_65;
  wire       [0:0]    _zz_sbuf_wdat_2_66;
  wire       [56:0]   _zz_sbuf_wdat_2_67;
  wire       [0:0]    _zz_sbuf_wdat_2_68;
  wire       [52:0]   _zz_sbuf_wdat_2_69;
  wire       [0:0]    _zz_sbuf_wdat_2_70;
  wire       [48:0]   _zz_sbuf_wdat_2_71;
  wire       [0:0]    _zz_sbuf_wdat_2_72;
  wire       [44:0]   _zz_sbuf_wdat_2_73;
  wire       [0:0]    _zz_sbuf_wdat_2_74;
  wire       [40:0]   _zz_sbuf_wdat_2_75;
  wire       [0:0]    _zz_sbuf_wdat_2_76;
  wire       [36:0]   _zz_sbuf_wdat_2_77;
  wire       [0:0]    _zz_sbuf_wdat_2_78;
  wire       [32:0]   _zz_sbuf_wdat_2_79;
  wire       [0:0]    _zz_sbuf_wdat_2_80;
  wire       [28:0]   _zz_sbuf_wdat_2_81;
  wire       [0:0]    _zz_sbuf_wdat_2_82;
  wire       [24:0]   _zz_sbuf_wdat_2_83;
  wire       [0:0]    _zz_sbuf_wdat_2_84;
  wire       [20:0]   _zz_sbuf_wdat_2_85;
  wire       [0:0]    _zz_sbuf_wdat_2_86;
  wire       [16:0]   _zz_sbuf_wdat_2_87;
  wire       [0:0]    _zz_sbuf_wdat_2_88;
  wire       [12:0]   _zz_sbuf_wdat_2_89;
  wire       [0:0]    _zz_sbuf_wdat_2_90;
  wire       [8:0]    _zz_sbuf_wdat_2_91;
  wire       [0:0]    _zz_sbuf_wdat_2_92;
  wire       [4:0]    _zz_sbuf_wdat_2_93;
  wire       [0:0]    _zz_sbuf_wdat_2_94;
  wire       [59:0]   _zz_sbuf_wdat_2_95;
  wire       [0:0]    _zz_sbuf_wdat_2_96;
  wire       [55:0]   _zz_sbuf_wdat_2_97;
  wire       [0:0]    _zz_sbuf_wdat_2_98;
  wire       [51:0]   _zz_sbuf_wdat_2_99;
  wire       [0:0]    _zz_sbuf_wdat_2_100;
  wire       [47:0]   _zz_sbuf_wdat_2_101;
  wire       [0:0]    _zz_sbuf_wdat_2_102;
  wire       [43:0]   _zz_sbuf_wdat_2_103;
  wire       [0:0]    _zz_sbuf_wdat_2_104;
  wire       [39:0]   _zz_sbuf_wdat_2_105;
  wire       [0:0]    _zz_sbuf_wdat_2_106;
  wire       [35:0]   _zz_sbuf_wdat_2_107;
  wire       [0:0]    _zz_sbuf_wdat_2_108;
  wire       [31:0]   _zz_sbuf_wdat_2_109;
  wire       [0:0]    _zz_sbuf_wdat_2_110;
  wire       [27:0]   _zz_sbuf_wdat_2_111;
  wire       [0:0]    _zz_sbuf_wdat_2_112;
  wire       [23:0]   _zz_sbuf_wdat_2_113;
  wire       [0:0]    _zz_sbuf_wdat_2_114;
  wire       [19:0]   _zz_sbuf_wdat_2_115;
  wire       [0:0]    _zz_sbuf_wdat_2_116;
  wire       [15:0]   _zz_sbuf_wdat_2_117;
  wire       [0:0]    _zz_sbuf_wdat_2_118;
  wire       [11:0]   _zz_sbuf_wdat_2_119;
  wire       [0:0]    _zz_sbuf_wdat_2_120;
  wire       [7:0]    _zz_sbuf_wdat_2_121;
  wire       [0:0]    _zz_sbuf_wdat_2_122;
  wire       [3:0]    _zz_sbuf_wdat_2_123;
  wire       [0:0]    _zz_sbuf_wdat_3;
  wire       [61:0]   _zz_sbuf_wdat_3_1;
  wire       [0:0]    _zz_sbuf_wdat_3_2;
  wire       [57:0]   _zz_sbuf_wdat_3_3;
  wire       [0:0]    _zz_sbuf_wdat_3_4;
  wire       [53:0]   _zz_sbuf_wdat_3_5;
  wire       [0:0]    _zz_sbuf_wdat_3_6;
  wire       [49:0]   _zz_sbuf_wdat_3_7;
  wire       [0:0]    _zz_sbuf_wdat_3_8;
  wire       [45:0]   _zz_sbuf_wdat_3_9;
  wire       [0:0]    _zz_sbuf_wdat_3_10;
  wire       [41:0]   _zz_sbuf_wdat_3_11;
  wire       [0:0]    _zz_sbuf_wdat_3_12;
  wire       [37:0]   _zz_sbuf_wdat_3_13;
  wire       [0:0]    _zz_sbuf_wdat_3_14;
  wire       [33:0]   _zz_sbuf_wdat_3_15;
  wire       [0:0]    _zz_sbuf_wdat_3_16;
  wire       [29:0]   _zz_sbuf_wdat_3_17;
  wire       [0:0]    _zz_sbuf_wdat_3_18;
  wire       [25:0]   _zz_sbuf_wdat_3_19;
  wire       [0:0]    _zz_sbuf_wdat_3_20;
  wire       [21:0]   _zz_sbuf_wdat_3_21;
  wire       [0:0]    _zz_sbuf_wdat_3_22;
  wire       [17:0]   _zz_sbuf_wdat_3_23;
  wire       [0:0]    _zz_sbuf_wdat_3_24;
  wire       [13:0]   _zz_sbuf_wdat_3_25;
  wire       [0:0]    _zz_sbuf_wdat_3_26;
  wire       [9:0]    _zz_sbuf_wdat_3_27;
  wire       [0:0]    _zz_sbuf_wdat_3_28;
  wire       [5:0]    _zz_sbuf_wdat_3_29;
  wire       [0:0]    _zz_sbuf_wdat_3_30;
  wire       [0:0]    _zz_sbuf_wdat_3_31;
  wire       [0:0]    _zz_sbuf_wdat_3_32;
  wire       [61:0]   _zz_sbuf_wdat_3_33;
  wire       [0:0]    _zz_sbuf_wdat_3_34;
  wire       [57:0]   _zz_sbuf_wdat_3_35;
  wire       [0:0]    _zz_sbuf_wdat_3_36;
  wire       [53:0]   _zz_sbuf_wdat_3_37;
  wire       [0:0]    _zz_sbuf_wdat_3_38;
  wire       [49:0]   _zz_sbuf_wdat_3_39;
  wire       [0:0]    _zz_sbuf_wdat_3_40;
  wire       [45:0]   _zz_sbuf_wdat_3_41;
  wire       [0:0]    _zz_sbuf_wdat_3_42;
  wire       [41:0]   _zz_sbuf_wdat_3_43;
  wire       [0:0]    _zz_sbuf_wdat_3_44;
  wire       [37:0]   _zz_sbuf_wdat_3_45;
  wire       [0:0]    _zz_sbuf_wdat_3_46;
  wire       [33:0]   _zz_sbuf_wdat_3_47;
  wire       [0:0]    _zz_sbuf_wdat_3_48;
  wire       [29:0]   _zz_sbuf_wdat_3_49;
  wire       [0:0]    _zz_sbuf_wdat_3_50;
  wire       [25:0]   _zz_sbuf_wdat_3_51;
  wire       [0:0]    _zz_sbuf_wdat_3_52;
  wire       [21:0]   _zz_sbuf_wdat_3_53;
  wire       [0:0]    _zz_sbuf_wdat_3_54;
  wire       [17:0]   _zz_sbuf_wdat_3_55;
  wire       [0:0]    _zz_sbuf_wdat_3_56;
  wire       [13:0]   _zz_sbuf_wdat_3_57;
  wire       [0:0]    _zz_sbuf_wdat_3_58;
  wire       [9:0]    _zz_sbuf_wdat_3_59;
  wire       [0:0]    _zz_sbuf_wdat_3_60;
  wire       [5:0]    _zz_sbuf_wdat_3_61;
  wire       [0:0]    _zz_sbuf_wdat_3_62;
  wire       [0:0]    _zz_sbuf_wdat_3_63;
  wire       [0:0]    _zz_sbuf_wdat_3_64;
  wire       [60:0]   _zz_sbuf_wdat_3_65;
  wire       [0:0]    _zz_sbuf_wdat_3_66;
  wire       [56:0]   _zz_sbuf_wdat_3_67;
  wire       [0:0]    _zz_sbuf_wdat_3_68;
  wire       [52:0]   _zz_sbuf_wdat_3_69;
  wire       [0:0]    _zz_sbuf_wdat_3_70;
  wire       [48:0]   _zz_sbuf_wdat_3_71;
  wire       [0:0]    _zz_sbuf_wdat_3_72;
  wire       [44:0]   _zz_sbuf_wdat_3_73;
  wire       [0:0]    _zz_sbuf_wdat_3_74;
  wire       [40:0]   _zz_sbuf_wdat_3_75;
  wire       [0:0]    _zz_sbuf_wdat_3_76;
  wire       [36:0]   _zz_sbuf_wdat_3_77;
  wire       [0:0]    _zz_sbuf_wdat_3_78;
  wire       [32:0]   _zz_sbuf_wdat_3_79;
  wire       [0:0]    _zz_sbuf_wdat_3_80;
  wire       [28:0]   _zz_sbuf_wdat_3_81;
  wire       [0:0]    _zz_sbuf_wdat_3_82;
  wire       [24:0]   _zz_sbuf_wdat_3_83;
  wire       [0:0]    _zz_sbuf_wdat_3_84;
  wire       [20:0]   _zz_sbuf_wdat_3_85;
  wire       [0:0]    _zz_sbuf_wdat_3_86;
  wire       [16:0]   _zz_sbuf_wdat_3_87;
  wire       [0:0]    _zz_sbuf_wdat_3_88;
  wire       [12:0]   _zz_sbuf_wdat_3_89;
  wire       [0:0]    _zz_sbuf_wdat_3_90;
  wire       [8:0]    _zz_sbuf_wdat_3_91;
  wire       [0:0]    _zz_sbuf_wdat_3_92;
  wire       [4:0]    _zz_sbuf_wdat_3_93;
  wire       [0:0]    _zz_sbuf_wdat_3_94;
  wire       [59:0]   _zz_sbuf_wdat_3_95;
  wire       [0:0]    _zz_sbuf_wdat_3_96;
  wire       [55:0]   _zz_sbuf_wdat_3_97;
  wire       [0:0]    _zz_sbuf_wdat_3_98;
  wire       [51:0]   _zz_sbuf_wdat_3_99;
  wire       [0:0]    _zz_sbuf_wdat_3_100;
  wire       [47:0]   _zz_sbuf_wdat_3_101;
  wire       [0:0]    _zz_sbuf_wdat_3_102;
  wire       [43:0]   _zz_sbuf_wdat_3_103;
  wire       [0:0]    _zz_sbuf_wdat_3_104;
  wire       [39:0]   _zz_sbuf_wdat_3_105;
  wire       [0:0]    _zz_sbuf_wdat_3_106;
  wire       [35:0]   _zz_sbuf_wdat_3_107;
  wire       [0:0]    _zz_sbuf_wdat_3_108;
  wire       [31:0]   _zz_sbuf_wdat_3_109;
  wire       [0:0]    _zz_sbuf_wdat_3_110;
  wire       [27:0]   _zz_sbuf_wdat_3_111;
  wire       [0:0]    _zz_sbuf_wdat_3_112;
  wire       [23:0]   _zz_sbuf_wdat_3_113;
  wire       [0:0]    _zz_sbuf_wdat_3_114;
  wire       [19:0]   _zz_sbuf_wdat_3_115;
  wire       [0:0]    _zz_sbuf_wdat_3_116;
  wire       [15:0]   _zz_sbuf_wdat_3_117;
  wire       [0:0]    _zz_sbuf_wdat_3_118;
  wire       [11:0]   _zz_sbuf_wdat_3_119;
  wire       [0:0]    _zz_sbuf_wdat_3_120;
  wire       [7:0]    _zz_sbuf_wdat_3_121;
  wire       [0:0]    _zz_sbuf_wdat_3_122;
  wire       [3:0]    _zz_sbuf_wdat_3_123;
  wire       [0:0]    _zz_sbuf_wdat_4;
  wire       [61:0]   _zz_sbuf_wdat_4_1;
  wire       [0:0]    _zz_sbuf_wdat_4_2;
  wire       [57:0]   _zz_sbuf_wdat_4_3;
  wire       [0:0]    _zz_sbuf_wdat_4_4;
  wire       [53:0]   _zz_sbuf_wdat_4_5;
  wire       [0:0]    _zz_sbuf_wdat_4_6;
  wire       [49:0]   _zz_sbuf_wdat_4_7;
  wire       [0:0]    _zz_sbuf_wdat_4_8;
  wire       [45:0]   _zz_sbuf_wdat_4_9;
  wire       [0:0]    _zz_sbuf_wdat_4_10;
  wire       [41:0]   _zz_sbuf_wdat_4_11;
  wire       [0:0]    _zz_sbuf_wdat_4_12;
  wire       [37:0]   _zz_sbuf_wdat_4_13;
  wire       [0:0]    _zz_sbuf_wdat_4_14;
  wire       [33:0]   _zz_sbuf_wdat_4_15;
  wire       [0:0]    _zz_sbuf_wdat_4_16;
  wire       [29:0]   _zz_sbuf_wdat_4_17;
  wire       [0:0]    _zz_sbuf_wdat_4_18;
  wire       [25:0]   _zz_sbuf_wdat_4_19;
  wire       [0:0]    _zz_sbuf_wdat_4_20;
  wire       [21:0]   _zz_sbuf_wdat_4_21;
  wire       [0:0]    _zz_sbuf_wdat_4_22;
  wire       [17:0]   _zz_sbuf_wdat_4_23;
  wire       [0:0]    _zz_sbuf_wdat_4_24;
  wire       [13:0]   _zz_sbuf_wdat_4_25;
  wire       [0:0]    _zz_sbuf_wdat_4_26;
  wire       [9:0]    _zz_sbuf_wdat_4_27;
  wire       [0:0]    _zz_sbuf_wdat_4_28;
  wire       [5:0]    _zz_sbuf_wdat_4_29;
  wire       [0:0]    _zz_sbuf_wdat_4_30;
  wire       [0:0]    _zz_sbuf_wdat_4_31;
  wire       [0:0]    _zz_sbuf_wdat_4_32;
  wire       [61:0]   _zz_sbuf_wdat_4_33;
  wire       [0:0]    _zz_sbuf_wdat_4_34;
  wire       [57:0]   _zz_sbuf_wdat_4_35;
  wire       [0:0]    _zz_sbuf_wdat_4_36;
  wire       [53:0]   _zz_sbuf_wdat_4_37;
  wire       [0:0]    _zz_sbuf_wdat_4_38;
  wire       [49:0]   _zz_sbuf_wdat_4_39;
  wire       [0:0]    _zz_sbuf_wdat_4_40;
  wire       [45:0]   _zz_sbuf_wdat_4_41;
  wire       [0:0]    _zz_sbuf_wdat_4_42;
  wire       [41:0]   _zz_sbuf_wdat_4_43;
  wire       [0:0]    _zz_sbuf_wdat_4_44;
  wire       [37:0]   _zz_sbuf_wdat_4_45;
  wire       [0:0]    _zz_sbuf_wdat_4_46;
  wire       [33:0]   _zz_sbuf_wdat_4_47;
  wire       [0:0]    _zz_sbuf_wdat_4_48;
  wire       [29:0]   _zz_sbuf_wdat_4_49;
  wire       [0:0]    _zz_sbuf_wdat_4_50;
  wire       [25:0]   _zz_sbuf_wdat_4_51;
  wire       [0:0]    _zz_sbuf_wdat_4_52;
  wire       [21:0]   _zz_sbuf_wdat_4_53;
  wire       [0:0]    _zz_sbuf_wdat_4_54;
  wire       [17:0]   _zz_sbuf_wdat_4_55;
  wire       [0:0]    _zz_sbuf_wdat_4_56;
  wire       [13:0]   _zz_sbuf_wdat_4_57;
  wire       [0:0]    _zz_sbuf_wdat_4_58;
  wire       [9:0]    _zz_sbuf_wdat_4_59;
  wire       [0:0]    _zz_sbuf_wdat_4_60;
  wire       [5:0]    _zz_sbuf_wdat_4_61;
  wire       [0:0]    _zz_sbuf_wdat_4_62;
  wire       [0:0]    _zz_sbuf_wdat_4_63;
  wire       [0:0]    _zz_sbuf_wdat_4_64;
  wire       [60:0]   _zz_sbuf_wdat_4_65;
  wire       [0:0]    _zz_sbuf_wdat_4_66;
  wire       [56:0]   _zz_sbuf_wdat_4_67;
  wire       [0:0]    _zz_sbuf_wdat_4_68;
  wire       [52:0]   _zz_sbuf_wdat_4_69;
  wire       [0:0]    _zz_sbuf_wdat_4_70;
  wire       [48:0]   _zz_sbuf_wdat_4_71;
  wire       [0:0]    _zz_sbuf_wdat_4_72;
  wire       [44:0]   _zz_sbuf_wdat_4_73;
  wire       [0:0]    _zz_sbuf_wdat_4_74;
  wire       [40:0]   _zz_sbuf_wdat_4_75;
  wire       [0:0]    _zz_sbuf_wdat_4_76;
  wire       [36:0]   _zz_sbuf_wdat_4_77;
  wire       [0:0]    _zz_sbuf_wdat_4_78;
  wire       [32:0]   _zz_sbuf_wdat_4_79;
  wire       [0:0]    _zz_sbuf_wdat_4_80;
  wire       [28:0]   _zz_sbuf_wdat_4_81;
  wire       [0:0]    _zz_sbuf_wdat_4_82;
  wire       [24:0]   _zz_sbuf_wdat_4_83;
  wire       [0:0]    _zz_sbuf_wdat_4_84;
  wire       [20:0]   _zz_sbuf_wdat_4_85;
  wire       [0:0]    _zz_sbuf_wdat_4_86;
  wire       [16:0]   _zz_sbuf_wdat_4_87;
  wire       [0:0]    _zz_sbuf_wdat_4_88;
  wire       [12:0]   _zz_sbuf_wdat_4_89;
  wire       [0:0]    _zz_sbuf_wdat_4_90;
  wire       [8:0]    _zz_sbuf_wdat_4_91;
  wire       [0:0]    _zz_sbuf_wdat_4_92;
  wire       [4:0]    _zz_sbuf_wdat_4_93;
  wire       [0:0]    _zz_sbuf_wdat_4_94;
  wire       [59:0]   _zz_sbuf_wdat_4_95;
  wire       [0:0]    _zz_sbuf_wdat_4_96;
  wire       [55:0]   _zz_sbuf_wdat_4_97;
  wire       [0:0]    _zz_sbuf_wdat_4_98;
  wire       [51:0]   _zz_sbuf_wdat_4_99;
  wire       [0:0]    _zz_sbuf_wdat_4_100;
  wire       [47:0]   _zz_sbuf_wdat_4_101;
  wire       [0:0]    _zz_sbuf_wdat_4_102;
  wire       [43:0]   _zz_sbuf_wdat_4_103;
  wire       [0:0]    _zz_sbuf_wdat_4_104;
  wire       [39:0]   _zz_sbuf_wdat_4_105;
  wire       [0:0]    _zz_sbuf_wdat_4_106;
  wire       [35:0]   _zz_sbuf_wdat_4_107;
  wire       [0:0]    _zz_sbuf_wdat_4_108;
  wire       [31:0]   _zz_sbuf_wdat_4_109;
  wire       [0:0]    _zz_sbuf_wdat_4_110;
  wire       [27:0]   _zz_sbuf_wdat_4_111;
  wire       [0:0]    _zz_sbuf_wdat_4_112;
  wire       [23:0]   _zz_sbuf_wdat_4_113;
  wire       [0:0]    _zz_sbuf_wdat_4_114;
  wire       [19:0]   _zz_sbuf_wdat_4_115;
  wire       [0:0]    _zz_sbuf_wdat_4_116;
  wire       [15:0]   _zz_sbuf_wdat_4_117;
  wire       [0:0]    _zz_sbuf_wdat_4_118;
  wire       [11:0]   _zz_sbuf_wdat_4_119;
  wire       [0:0]    _zz_sbuf_wdat_4_120;
  wire       [7:0]    _zz_sbuf_wdat_4_121;
  wire       [0:0]    _zz_sbuf_wdat_4_122;
  wire       [3:0]    _zz_sbuf_wdat_4_123;
  wire       [0:0]    _zz_sbuf_wdat_5;
  wire       [61:0]   _zz_sbuf_wdat_5_1;
  wire       [0:0]    _zz_sbuf_wdat_5_2;
  wire       [57:0]   _zz_sbuf_wdat_5_3;
  wire       [0:0]    _zz_sbuf_wdat_5_4;
  wire       [53:0]   _zz_sbuf_wdat_5_5;
  wire       [0:0]    _zz_sbuf_wdat_5_6;
  wire       [49:0]   _zz_sbuf_wdat_5_7;
  wire       [0:0]    _zz_sbuf_wdat_5_8;
  wire       [45:0]   _zz_sbuf_wdat_5_9;
  wire       [0:0]    _zz_sbuf_wdat_5_10;
  wire       [41:0]   _zz_sbuf_wdat_5_11;
  wire       [0:0]    _zz_sbuf_wdat_5_12;
  wire       [37:0]   _zz_sbuf_wdat_5_13;
  wire       [0:0]    _zz_sbuf_wdat_5_14;
  wire       [33:0]   _zz_sbuf_wdat_5_15;
  wire       [0:0]    _zz_sbuf_wdat_5_16;
  wire       [29:0]   _zz_sbuf_wdat_5_17;
  wire       [0:0]    _zz_sbuf_wdat_5_18;
  wire       [25:0]   _zz_sbuf_wdat_5_19;
  wire       [0:0]    _zz_sbuf_wdat_5_20;
  wire       [21:0]   _zz_sbuf_wdat_5_21;
  wire       [0:0]    _zz_sbuf_wdat_5_22;
  wire       [17:0]   _zz_sbuf_wdat_5_23;
  wire       [0:0]    _zz_sbuf_wdat_5_24;
  wire       [13:0]   _zz_sbuf_wdat_5_25;
  wire       [0:0]    _zz_sbuf_wdat_5_26;
  wire       [9:0]    _zz_sbuf_wdat_5_27;
  wire       [0:0]    _zz_sbuf_wdat_5_28;
  wire       [5:0]    _zz_sbuf_wdat_5_29;
  wire       [0:0]    _zz_sbuf_wdat_5_30;
  wire       [0:0]    _zz_sbuf_wdat_5_31;
  wire       [0:0]    _zz_sbuf_wdat_5_32;
  wire       [61:0]   _zz_sbuf_wdat_5_33;
  wire       [0:0]    _zz_sbuf_wdat_5_34;
  wire       [57:0]   _zz_sbuf_wdat_5_35;
  wire       [0:0]    _zz_sbuf_wdat_5_36;
  wire       [53:0]   _zz_sbuf_wdat_5_37;
  wire       [0:0]    _zz_sbuf_wdat_5_38;
  wire       [49:0]   _zz_sbuf_wdat_5_39;
  wire       [0:0]    _zz_sbuf_wdat_5_40;
  wire       [45:0]   _zz_sbuf_wdat_5_41;
  wire       [0:0]    _zz_sbuf_wdat_5_42;
  wire       [41:0]   _zz_sbuf_wdat_5_43;
  wire       [0:0]    _zz_sbuf_wdat_5_44;
  wire       [37:0]   _zz_sbuf_wdat_5_45;
  wire       [0:0]    _zz_sbuf_wdat_5_46;
  wire       [33:0]   _zz_sbuf_wdat_5_47;
  wire       [0:0]    _zz_sbuf_wdat_5_48;
  wire       [29:0]   _zz_sbuf_wdat_5_49;
  wire       [0:0]    _zz_sbuf_wdat_5_50;
  wire       [25:0]   _zz_sbuf_wdat_5_51;
  wire       [0:0]    _zz_sbuf_wdat_5_52;
  wire       [21:0]   _zz_sbuf_wdat_5_53;
  wire       [0:0]    _zz_sbuf_wdat_5_54;
  wire       [17:0]   _zz_sbuf_wdat_5_55;
  wire       [0:0]    _zz_sbuf_wdat_5_56;
  wire       [13:0]   _zz_sbuf_wdat_5_57;
  wire       [0:0]    _zz_sbuf_wdat_5_58;
  wire       [9:0]    _zz_sbuf_wdat_5_59;
  wire       [0:0]    _zz_sbuf_wdat_5_60;
  wire       [5:0]    _zz_sbuf_wdat_5_61;
  wire       [0:0]    _zz_sbuf_wdat_5_62;
  wire       [0:0]    _zz_sbuf_wdat_5_63;
  wire       [0:0]    _zz_sbuf_wdat_5_64;
  wire       [60:0]   _zz_sbuf_wdat_5_65;
  wire       [0:0]    _zz_sbuf_wdat_5_66;
  wire       [56:0]   _zz_sbuf_wdat_5_67;
  wire       [0:0]    _zz_sbuf_wdat_5_68;
  wire       [52:0]   _zz_sbuf_wdat_5_69;
  wire       [0:0]    _zz_sbuf_wdat_5_70;
  wire       [48:0]   _zz_sbuf_wdat_5_71;
  wire       [0:0]    _zz_sbuf_wdat_5_72;
  wire       [44:0]   _zz_sbuf_wdat_5_73;
  wire       [0:0]    _zz_sbuf_wdat_5_74;
  wire       [40:0]   _zz_sbuf_wdat_5_75;
  wire       [0:0]    _zz_sbuf_wdat_5_76;
  wire       [36:0]   _zz_sbuf_wdat_5_77;
  wire       [0:0]    _zz_sbuf_wdat_5_78;
  wire       [32:0]   _zz_sbuf_wdat_5_79;
  wire       [0:0]    _zz_sbuf_wdat_5_80;
  wire       [28:0]   _zz_sbuf_wdat_5_81;
  wire       [0:0]    _zz_sbuf_wdat_5_82;
  wire       [24:0]   _zz_sbuf_wdat_5_83;
  wire       [0:0]    _zz_sbuf_wdat_5_84;
  wire       [20:0]   _zz_sbuf_wdat_5_85;
  wire       [0:0]    _zz_sbuf_wdat_5_86;
  wire       [16:0]   _zz_sbuf_wdat_5_87;
  wire       [0:0]    _zz_sbuf_wdat_5_88;
  wire       [12:0]   _zz_sbuf_wdat_5_89;
  wire       [0:0]    _zz_sbuf_wdat_5_90;
  wire       [8:0]    _zz_sbuf_wdat_5_91;
  wire       [0:0]    _zz_sbuf_wdat_5_92;
  wire       [4:0]    _zz_sbuf_wdat_5_93;
  wire       [0:0]    _zz_sbuf_wdat_5_94;
  wire       [59:0]   _zz_sbuf_wdat_5_95;
  wire       [0:0]    _zz_sbuf_wdat_5_96;
  wire       [55:0]   _zz_sbuf_wdat_5_97;
  wire       [0:0]    _zz_sbuf_wdat_5_98;
  wire       [51:0]   _zz_sbuf_wdat_5_99;
  wire       [0:0]    _zz_sbuf_wdat_5_100;
  wire       [47:0]   _zz_sbuf_wdat_5_101;
  wire       [0:0]    _zz_sbuf_wdat_5_102;
  wire       [43:0]   _zz_sbuf_wdat_5_103;
  wire       [0:0]    _zz_sbuf_wdat_5_104;
  wire       [39:0]   _zz_sbuf_wdat_5_105;
  wire       [0:0]    _zz_sbuf_wdat_5_106;
  wire       [35:0]   _zz_sbuf_wdat_5_107;
  wire       [0:0]    _zz_sbuf_wdat_5_108;
  wire       [31:0]   _zz_sbuf_wdat_5_109;
  wire       [0:0]    _zz_sbuf_wdat_5_110;
  wire       [27:0]   _zz_sbuf_wdat_5_111;
  wire       [0:0]    _zz_sbuf_wdat_5_112;
  wire       [23:0]   _zz_sbuf_wdat_5_113;
  wire       [0:0]    _zz_sbuf_wdat_5_114;
  wire       [19:0]   _zz_sbuf_wdat_5_115;
  wire       [0:0]    _zz_sbuf_wdat_5_116;
  wire       [15:0]   _zz_sbuf_wdat_5_117;
  wire       [0:0]    _zz_sbuf_wdat_5_118;
  wire       [11:0]   _zz_sbuf_wdat_5_119;
  wire       [0:0]    _zz_sbuf_wdat_5_120;
  wire       [7:0]    _zz_sbuf_wdat_5_121;
  wire       [0:0]    _zz_sbuf_wdat_5_122;
  wire       [3:0]    _zz_sbuf_wdat_5_123;
  wire       [0:0]    _zz_sbuf_wdat_6;
  wire       [61:0]   _zz_sbuf_wdat_6_1;
  wire       [0:0]    _zz_sbuf_wdat_6_2;
  wire       [57:0]   _zz_sbuf_wdat_6_3;
  wire       [0:0]    _zz_sbuf_wdat_6_4;
  wire       [53:0]   _zz_sbuf_wdat_6_5;
  wire       [0:0]    _zz_sbuf_wdat_6_6;
  wire       [49:0]   _zz_sbuf_wdat_6_7;
  wire       [0:0]    _zz_sbuf_wdat_6_8;
  wire       [45:0]   _zz_sbuf_wdat_6_9;
  wire       [0:0]    _zz_sbuf_wdat_6_10;
  wire       [41:0]   _zz_sbuf_wdat_6_11;
  wire       [0:0]    _zz_sbuf_wdat_6_12;
  wire       [37:0]   _zz_sbuf_wdat_6_13;
  wire       [0:0]    _zz_sbuf_wdat_6_14;
  wire       [33:0]   _zz_sbuf_wdat_6_15;
  wire       [0:0]    _zz_sbuf_wdat_6_16;
  wire       [29:0]   _zz_sbuf_wdat_6_17;
  wire       [0:0]    _zz_sbuf_wdat_6_18;
  wire       [25:0]   _zz_sbuf_wdat_6_19;
  wire       [0:0]    _zz_sbuf_wdat_6_20;
  wire       [21:0]   _zz_sbuf_wdat_6_21;
  wire       [0:0]    _zz_sbuf_wdat_6_22;
  wire       [17:0]   _zz_sbuf_wdat_6_23;
  wire       [0:0]    _zz_sbuf_wdat_6_24;
  wire       [13:0]   _zz_sbuf_wdat_6_25;
  wire       [0:0]    _zz_sbuf_wdat_6_26;
  wire       [9:0]    _zz_sbuf_wdat_6_27;
  wire       [0:0]    _zz_sbuf_wdat_6_28;
  wire       [5:0]    _zz_sbuf_wdat_6_29;
  wire       [0:0]    _zz_sbuf_wdat_6_30;
  wire       [0:0]    _zz_sbuf_wdat_6_31;
  wire       [0:0]    _zz_sbuf_wdat_6_32;
  wire       [61:0]   _zz_sbuf_wdat_6_33;
  wire       [0:0]    _zz_sbuf_wdat_6_34;
  wire       [57:0]   _zz_sbuf_wdat_6_35;
  wire       [0:0]    _zz_sbuf_wdat_6_36;
  wire       [53:0]   _zz_sbuf_wdat_6_37;
  wire       [0:0]    _zz_sbuf_wdat_6_38;
  wire       [49:0]   _zz_sbuf_wdat_6_39;
  wire       [0:0]    _zz_sbuf_wdat_6_40;
  wire       [45:0]   _zz_sbuf_wdat_6_41;
  wire       [0:0]    _zz_sbuf_wdat_6_42;
  wire       [41:0]   _zz_sbuf_wdat_6_43;
  wire       [0:0]    _zz_sbuf_wdat_6_44;
  wire       [37:0]   _zz_sbuf_wdat_6_45;
  wire       [0:0]    _zz_sbuf_wdat_6_46;
  wire       [33:0]   _zz_sbuf_wdat_6_47;
  wire       [0:0]    _zz_sbuf_wdat_6_48;
  wire       [29:0]   _zz_sbuf_wdat_6_49;
  wire       [0:0]    _zz_sbuf_wdat_6_50;
  wire       [25:0]   _zz_sbuf_wdat_6_51;
  wire       [0:0]    _zz_sbuf_wdat_6_52;
  wire       [21:0]   _zz_sbuf_wdat_6_53;
  wire       [0:0]    _zz_sbuf_wdat_6_54;
  wire       [17:0]   _zz_sbuf_wdat_6_55;
  wire       [0:0]    _zz_sbuf_wdat_6_56;
  wire       [13:0]   _zz_sbuf_wdat_6_57;
  wire       [0:0]    _zz_sbuf_wdat_6_58;
  wire       [9:0]    _zz_sbuf_wdat_6_59;
  wire       [0:0]    _zz_sbuf_wdat_6_60;
  wire       [5:0]    _zz_sbuf_wdat_6_61;
  wire       [0:0]    _zz_sbuf_wdat_6_62;
  wire       [0:0]    _zz_sbuf_wdat_6_63;
  wire       [0:0]    _zz_sbuf_wdat_6_64;
  wire       [60:0]   _zz_sbuf_wdat_6_65;
  wire       [0:0]    _zz_sbuf_wdat_6_66;
  wire       [56:0]   _zz_sbuf_wdat_6_67;
  wire       [0:0]    _zz_sbuf_wdat_6_68;
  wire       [52:0]   _zz_sbuf_wdat_6_69;
  wire       [0:0]    _zz_sbuf_wdat_6_70;
  wire       [48:0]   _zz_sbuf_wdat_6_71;
  wire       [0:0]    _zz_sbuf_wdat_6_72;
  wire       [44:0]   _zz_sbuf_wdat_6_73;
  wire       [0:0]    _zz_sbuf_wdat_6_74;
  wire       [40:0]   _zz_sbuf_wdat_6_75;
  wire       [0:0]    _zz_sbuf_wdat_6_76;
  wire       [36:0]   _zz_sbuf_wdat_6_77;
  wire       [0:0]    _zz_sbuf_wdat_6_78;
  wire       [32:0]   _zz_sbuf_wdat_6_79;
  wire       [0:0]    _zz_sbuf_wdat_6_80;
  wire       [28:0]   _zz_sbuf_wdat_6_81;
  wire       [0:0]    _zz_sbuf_wdat_6_82;
  wire       [24:0]   _zz_sbuf_wdat_6_83;
  wire       [0:0]    _zz_sbuf_wdat_6_84;
  wire       [20:0]   _zz_sbuf_wdat_6_85;
  wire       [0:0]    _zz_sbuf_wdat_6_86;
  wire       [16:0]   _zz_sbuf_wdat_6_87;
  wire       [0:0]    _zz_sbuf_wdat_6_88;
  wire       [12:0]   _zz_sbuf_wdat_6_89;
  wire       [0:0]    _zz_sbuf_wdat_6_90;
  wire       [8:0]    _zz_sbuf_wdat_6_91;
  wire       [0:0]    _zz_sbuf_wdat_6_92;
  wire       [4:0]    _zz_sbuf_wdat_6_93;
  wire       [0:0]    _zz_sbuf_wdat_6_94;
  wire       [59:0]   _zz_sbuf_wdat_6_95;
  wire       [0:0]    _zz_sbuf_wdat_6_96;
  wire       [55:0]   _zz_sbuf_wdat_6_97;
  wire       [0:0]    _zz_sbuf_wdat_6_98;
  wire       [51:0]   _zz_sbuf_wdat_6_99;
  wire       [0:0]    _zz_sbuf_wdat_6_100;
  wire       [47:0]   _zz_sbuf_wdat_6_101;
  wire       [0:0]    _zz_sbuf_wdat_6_102;
  wire       [43:0]   _zz_sbuf_wdat_6_103;
  wire       [0:0]    _zz_sbuf_wdat_6_104;
  wire       [39:0]   _zz_sbuf_wdat_6_105;
  wire       [0:0]    _zz_sbuf_wdat_6_106;
  wire       [35:0]   _zz_sbuf_wdat_6_107;
  wire       [0:0]    _zz_sbuf_wdat_6_108;
  wire       [31:0]   _zz_sbuf_wdat_6_109;
  wire       [0:0]    _zz_sbuf_wdat_6_110;
  wire       [27:0]   _zz_sbuf_wdat_6_111;
  wire       [0:0]    _zz_sbuf_wdat_6_112;
  wire       [23:0]   _zz_sbuf_wdat_6_113;
  wire       [0:0]    _zz_sbuf_wdat_6_114;
  wire       [19:0]   _zz_sbuf_wdat_6_115;
  wire       [0:0]    _zz_sbuf_wdat_6_116;
  wire       [15:0]   _zz_sbuf_wdat_6_117;
  wire       [0:0]    _zz_sbuf_wdat_6_118;
  wire       [11:0]   _zz_sbuf_wdat_6_119;
  wire       [0:0]    _zz_sbuf_wdat_6_120;
  wire       [7:0]    _zz_sbuf_wdat_6_121;
  wire       [0:0]    _zz_sbuf_wdat_6_122;
  wire       [3:0]    _zz_sbuf_wdat_6_123;
  wire       [0:0]    _zz_sbuf_wdat_7;
  wire       [61:0]   _zz_sbuf_wdat_7_1;
  wire       [0:0]    _zz_sbuf_wdat_7_2;
  wire       [57:0]   _zz_sbuf_wdat_7_3;
  wire       [0:0]    _zz_sbuf_wdat_7_4;
  wire       [53:0]   _zz_sbuf_wdat_7_5;
  wire       [0:0]    _zz_sbuf_wdat_7_6;
  wire       [49:0]   _zz_sbuf_wdat_7_7;
  wire       [0:0]    _zz_sbuf_wdat_7_8;
  wire       [45:0]   _zz_sbuf_wdat_7_9;
  wire       [0:0]    _zz_sbuf_wdat_7_10;
  wire       [41:0]   _zz_sbuf_wdat_7_11;
  wire       [0:0]    _zz_sbuf_wdat_7_12;
  wire       [37:0]   _zz_sbuf_wdat_7_13;
  wire       [0:0]    _zz_sbuf_wdat_7_14;
  wire       [33:0]   _zz_sbuf_wdat_7_15;
  wire       [0:0]    _zz_sbuf_wdat_7_16;
  wire       [29:0]   _zz_sbuf_wdat_7_17;
  wire       [0:0]    _zz_sbuf_wdat_7_18;
  wire       [25:0]   _zz_sbuf_wdat_7_19;
  wire       [0:0]    _zz_sbuf_wdat_7_20;
  wire       [21:0]   _zz_sbuf_wdat_7_21;
  wire       [0:0]    _zz_sbuf_wdat_7_22;
  wire       [17:0]   _zz_sbuf_wdat_7_23;
  wire       [0:0]    _zz_sbuf_wdat_7_24;
  wire       [13:0]   _zz_sbuf_wdat_7_25;
  wire       [0:0]    _zz_sbuf_wdat_7_26;
  wire       [9:0]    _zz_sbuf_wdat_7_27;
  wire       [0:0]    _zz_sbuf_wdat_7_28;
  wire       [5:0]    _zz_sbuf_wdat_7_29;
  wire       [0:0]    _zz_sbuf_wdat_7_30;
  wire       [0:0]    _zz_sbuf_wdat_7_31;
  wire       [0:0]    _zz_sbuf_wdat_7_32;
  wire       [61:0]   _zz_sbuf_wdat_7_33;
  wire       [0:0]    _zz_sbuf_wdat_7_34;
  wire       [57:0]   _zz_sbuf_wdat_7_35;
  wire       [0:0]    _zz_sbuf_wdat_7_36;
  wire       [53:0]   _zz_sbuf_wdat_7_37;
  wire       [0:0]    _zz_sbuf_wdat_7_38;
  wire       [49:0]   _zz_sbuf_wdat_7_39;
  wire       [0:0]    _zz_sbuf_wdat_7_40;
  wire       [45:0]   _zz_sbuf_wdat_7_41;
  wire       [0:0]    _zz_sbuf_wdat_7_42;
  wire       [41:0]   _zz_sbuf_wdat_7_43;
  wire       [0:0]    _zz_sbuf_wdat_7_44;
  wire       [37:0]   _zz_sbuf_wdat_7_45;
  wire       [0:0]    _zz_sbuf_wdat_7_46;
  wire       [33:0]   _zz_sbuf_wdat_7_47;
  wire       [0:0]    _zz_sbuf_wdat_7_48;
  wire       [29:0]   _zz_sbuf_wdat_7_49;
  wire       [0:0]    _zz_sbuf_wdat_7_50;
  wire       [25:0]   _zz_sbuf_wdat_7_51;
  wire       [0:0]    _zz_sbuf_wdat_7_52;
  wire       [21:0]   _zz_sbuf_wdat_7_53;
  wire       [0:0]    _zz_sbuf_wdat_7_54;
  wire       [17:0]   _zz_sbuf_wdat_7_55;
  wire       [0:0]    _zz_sbuf_wdat_7_56;
  wire       [13:0]   _zz_sbuf_wdat_7_57;
  wire       [0:0]    _zz_sbuf_wdat_7_58;
  wire       [9:0]    _zz_sbuf_wdat_7_59;
  wire       [0:0]    _zz_sbuf_wdat_7_60;
  wire       [5:0]    _zz_sbuf_wdat_7_61;
  wire       [0:0]    _zz_sbuf_wdat_7_62;
  wire       [0:0]    _zz_sbuf_wdat_7_63;
  wire       [0:0]    _zz_sbuf_wdat_7_64;
  wire       [60:0]   _zz_sbuf_wdat_7_65;
  wire       [0:0]    _zz_sbuf_wdat_7_66;
  wire       [56:0]   _zz_sbuf_wdat_7_67;
  wire       [0:0]    _zz_sbuf_wdat_7_68;
  wire       [52:0]   _zz_sbuf_wdat_7_69;
  wire       [0:0]    _zz_sbuf_wdat_7_70;
  wire       [48:0]   _zz_sbuf_wdat_7_71;
  wire       [0:0]    _zz_sbuf_wdat_7_72;
  wire       [44:0]   _zz_sbuf_wdat_7_73;
  wire       [0:0]    _zz_sbuf_wdat_7_74;
  wire       [40:0]   _zz_sbuf_wdat_7_75;
  wire       [0:0]    _zz_sbuf_wdat_7_76;
  wire       [36:0]   _zz_sbuf_wdat_7_77;
  wire       [0:0]    _zz_sbuf_wdat_7_78;
  wire       [32:0]   _zz_sbuf_wdat_7_79;
  wire       [0:0]    _zz_sbuf_wdat_7_80;
  wire       [28:0]   _zz_sbuf_wdat_7_81;
  wire       [0:0]    _zz_sbuf_wdat_7_82;
  wire       [24:0]   _zz_sbuf_wdat_7_83;
  wire       [0:0]    _zz_sbuf_wdat_7_84;
  wire       [20:0]   _zz_sbuf_wdat_7_85;
  wire       [0:0]    _zz_sbuf_wdat_7_86;
  wire       [16:0]   _zz_sbuf_wdat_7_87;
  wire       [0:0]    _zz_sbuf_wdat_7_88;
  wire       [12:0]   _zz_sbuf_wdat_7_89;
  wire       [0:0]    _zz_sbuf_wdat_7_90;
  wire       [8:0]    _zz_sbuf_wdat_7_91;
  wire       [0:0]    _zz_sbuf_wdat_7_92;
  wire       [4:0]    _zz_sbuf_wdat_7_93;
  wire       [0:0]    _zz_sbuf_wdat_7_94;
  wire       [59:0]   _zz_sbuf_wdat_7_95;
  wire       [0:0]    _zz_sbuf_wdat_7_96;
  wire       [55:0]   _zz_sbuf_wdat_7_97;
  wire       [0:0]    _zz_sbuf_wdat_7_98;
  wire       [51:0]   _zz_sbuf_wdat_7_99;
  wire       [0:0]    _zz_sbuf_wdat_7_100;
  wire       [47:0]   _zz_sbuf_wdat_7_101;
  wire       [0:0]    _zz_sbuf_wdat_7_102;
  wire       [43:0]   _zz_sbuf_wdat_7_103;
  wire       [0:0]    _zz_sbuf_wdat_7_104;
  wire       [39:0]   _zz_sbuf_wdat_7_105;
  wire       [0:0]    _zz_sbuf_wdat_7_106;
  wire       [35:0]   _zz_sbuf_wdat_7_107;
  wire       [0:0]    _zz_sbuf_wdat_7_108;
  wire       [31:0]   _zz_sbuf_wdat_7_109;
  wire       [0:0]    _zz_sbuf_wdat_7_110;
  wire       [27:0]   _zz_sbuf_wdat_7_111;
  wire       [0:0]    _zz_sbuf_wdat_7_112;
  wire       [23:0]   _zz_sbuf_wdat_7_113;
  wire       [0:0]    _zz_sbuf_wdat_7_114;
  wire       [19:0]   _zz_sbuf_wdat_7_115;
  wire       [0:0]    _zz_sbuf_wdat_7_116;
  wire       [15:0]   _zz_sbuf_wdat_7_117;
  wire       [0:0]    _zz_sbuf_wdat_7_118;
  wire       [11:0]   _zz_sbuf_wdat_7_119;
  wire       [0:0]    _zz_sbuf_wdat_7_120;
  wire       [7:0]    _zz_sbuf_wdat_7_121;
  wire       [0:0]    _zz_sbuf_wdat_7_122;
  wire       [3:0]    _zz_sbuf_wdat_7_123;
  wire       [0:0]    _zz_sbuf_wdat_8;
  wire       [61:0]   _zz_sbuf_wdat_8_1;
  wire       [0:0]    _zz_sbuf_wdat_8_2;
  wire       [57:0]   _zz_sbuf_wdat_8_3;
  wire       [0:0]    _zz_sbuf_wdat_8_4;
  wire       [53:0]   _zz_sbuf_wdat_8_5;
  wire       [0:0]    _zz_sbuf_wdat_8_6;
  wire       [49:0]   _zz_sbuf_wdat_8_7;
  wire       [0:0]    _zz_sbuf_wdat_8_8;
  wire       [45:0]   _zz_sbuf_wdat_8_9;
  wire       [0:0]    _zz_sbuf_wdat_8_10;
  wire       [41:0]   _zz_sbuf_wdat_8_11;
  wire       [0:0]    _zz_sbuf_wdat_8_12;
  wire       [37:0]   _zz_sbuf_wdat_8_13;
  wire       [0:0]    _zz_sbuf_wdat_8_14;
  wire       [33:0]   _zz_sbuf_wdat_8_15;
  wire       [0:0]    _zz_sbuf_wdat_8_16;
  wire       [29:0]   _zz_sbuf_wdat_8_17;
  wire       [0:0]    _zz_sbuf_wdat_8_18;
  wire       [25:0]   _zz_sbuf_wdat_8_19;
  wire       [0:0]    _zz_sbuf_wdat_8_20;
  wire       [21:0]   _zz_sbuf_wdat_8_21;
  wire       [0:0]    _zz_sbuf_wdat_8_22;
  wire       [17:0]   _zz_sbuf_wdat_8_23;
  wire       [0:0]    _zz_sbuf_wdat_8_24;
  wire       [13:0]   _zz_sbuf_wdat_8_25;
  wire       [0:0]    _zz_sbuf_wdat_8_26;
  wire       [9:0]    _zz_sbuf_wdat_8_27;
  wire       [0:0]    _zz_sbuf_wdat_8_28;
  wire       [5:0]    _zz_sbuf_wdat_8_29;
  wire       [0:0]    _zz_sbuf_wdat_8_30;
  wire       [0:0]    _zz_sbuf_wdat_8_31;
  wire       [0:0]    _zz_sbuf_wdat_8_32;
  wire       [61:0]   _zz_sbuf_wdat_8_33;
  wire       [0:0]    _zz_sbuf_wdat_8_34;
  wire       [57:0]   _zz_sbuf_wdat_8_35;
  wire       [0:0]    _zz_sbuf_wdat_8_36;
  wire       [53:0]   _zz_sbuf_wdat_8_37;
  wire       [0:0]    _zz_sbuf_wdat_8_38;
  wire       [49:0]   _zz_sbuf_wdat_8_39;
  wire       [0:0]    _zz_sbuf_wdat_8_40;
  wire       [45:0]   _zz_sbuf_wdat_8_41;
  wire       [0:0]    _zz_sbuf_wdat_8_42;
  wire       [41:0]   _zz_sbuf_wdat_8_43;
  wire       [0:0]    _zz_sbuf_wdat_8_44;
  wire       [37:0]   _zz_sbuf_wdat_8_45;
  wire       [0:0]    _zz_sbuf_wdat_8_46;
  wire       [33:0]   _zz_sbuf_wdat_8_47;
  wire       [0:0]    _zz_sbuf_wdat_8_48;
  wire       [29:0]   _zz_sbuf_wdat_8_49;
  wire       [0:0]    _zz_sbuf_wdat_8_50;
  wire       [25:0]   _zz_sbuf_wdat_8_51;
  wire       [0:0]    _zz_sbuf_wdat_8_52;
  wire       [21:0]   _zz_sbuf_wdat_8_53;
  wire       [0:0]    _zz_sbuf_wdat_8_54;
  wire       [17:0]   _zz_sbuf_wdat_8_55;
  wire       [0:0]    _zz_sbuf_wdat_8_56;
  wire       [13:0]   _zz_sbuf_wdat_8_57;
  wire       [0:0]    _zz_sbuf_wdat_8_58;
  wire       [9:0]    _zz_sbuf_wdat_8_59;
  wire       [0:0]    _zz_sbuf_wdat_8_60;
  wire       [5:0]    _zz_sbuf_wdat_8_61;
  wire       [0:0]    _zz_sbuf_wdat_8_62;
  wire       [0:0]    _zz_sbuf_wdat_8_63;
  wire       [0:0]    _zz_sbuf_wdat_8_64;
  wire       [60:0]   _zz_sbuf_wdat_8_65;
  wire       [0:0]    _zz_sbuf_wdat_8_66;
  wire       [56:0]   _zz_sbuf_wdat_8_67;
  wire       [0:0]    _zz_sbuf_wdat_8_68;
  wire       [52:0]   _zz_sbuf_wdat_8_69;
  wire       [0:0]    _zz_sbuf_wdat_8_70;
  wire       [48:0]   _zz_sbuf_wdat_8_71;
  wire       [0:0]    _zz_sbuf_wdat_8_72;
  wire       [44:0]   _zz_sbuf_wdat_8_73;
  wire       [0:0]    _zz_sbuf_wdat_8_74;
  wire       [40:0]   _zz_sbuf_wdat_8_75;
  wire       [0:0]    _zz_sbuf_wdat_8_76;
  wire       [36:0]   _zz_sbuf_wdat_8_77;
  wire       [0:0]    _zz_sbuf_wdat_8_78;
  wire       [32:0]   _zz_sbuf_wdat_8_79;
  wire       [0:0]    _zz_sbuf_wdat_8_80;
  wire       [28:0]   _zz_sbuf_wdat_8_81;
  wire       [0:0]    _zz_sbuf_wdat_8_82;
  wire       [24:0]   _zz_sbuf_wdat_8_83;
  wire       [0:0]    _zz_sbuf_wdat_8_84;
  wire       [20:0]   _zz_sbuf_wdat_8_85;
  wire       [0:0]    _zz_sbuf_wdat_8_86;
  wire       [16:0]   _zz_sbuf_wdat_8_87;
  wire       [0:0]    _zz_sbuf_wdat_8_88;
  wire       [12:0]   _zz_sbuf_wdat_8_89;
  wire       [0:0]    _zz_sbuf_wdat_8_90;
  wire       [8:0]    _zz_sbuf_wdat_8_91;
  wire       [0:0]    _zz_sbuf_wdat_8_92;
  wire       [4:0]    _zz_sbuf_wdat_8_93;
  wire       [0:0]    _zz_sbuf_wdat_8_94;
  wire       [59:0]   _zz_sbuf_wdat_8_95;
  wire       [0:0]    _zz_sbuf_wdat_8_96;
  wire       [55:0]   _zz_sbuf_wdat_8_97;
  wire       [0:0]    _zz_sbuf_wdat_8_98;
  wire       [51:0]   _zz_sbuf_wdat_8_99;
  wire       [0:0]    _zz_sbuf_wdat_8_100;
  wire       [47:0]   _zz_sbuf_wdat_8_101;
  wire       [0:0]    _zz_sbuf_wdat_8_102;
  wire       [43:0]   _zz_sbuf_wdat_8_103;
  wire       [0:0]    _zz_sbuf_wdat_8_104;
  wire       [39:0]   _zz_sbuf_wdat_8_105;
  wire       [0:0]    _zz_sbuf_wdat_8_106;
  wire       [35:0]   _zz_sbuf_wdat_8_107;
  wire       [0:0]    _zz_sbuf_wdat_8_108;
  wire       [31:0]   _zz_sbuf_wdat_8_109;
  wire       [0:0]    _zz_sbuf_wdat_8_110;
  wire       [27:0]   _zz_sbuf_wdat_8_111;
  wire       [0:0]    _zz_sbuf_wdat_8_112;
  wire       [23:0]   _zz_sbuf_wdat_8_113;
  wire       [0:0]    _zz_sbuf_wdat_8_114;
  wire       [19:0]   _zz_sbuf_wdat_8_115;
  wire       [0:0]    _zz_sbuf_wdat_8_116;
  wire       [15:0]   _zz_sbuf_wdat_8_117;
  wire       [0:0]    _zz_sbuf_wdat_8_118;
  wire       [11:0]   _zz_sbuf_wdat_8_119;
  wire       [0:0]    _zz_sbuf_wdat_8_120;
  wire       [7:0]    _zz_sbuf_wdat_8_121;
  wire       [0:0]    _zz_sbuf_wdat_8_122;
  wire       [3:0]    _zz_sbuf_wdat_8_123;
  wire       [0:0]    _zz_sbuf_wdat_9;
  wire       [61:0]   _zz_sbuf_wdat_9_1;
  wire       [0:0]    _zz_sbuf_wdat_9_2;
  wire       [57:0]   _zz_sbuf_wdat_9_3;
  wire       [0:0]    _zz_sbuf_wdat_9_4;
  wire       [53:0]   _zz_sbuf_wdat_9_5;
  wire       [0:0]    _zz_sbuf_wdat_9_6;
  wire       [49:0]   _zz_sbuf_wdat_9_7;
  wire       [0:0]    _zz_sbuf_wdat_9_8;
  wire       [45:0]   _zz_sbuf_wdat_9_9;
  wire       [0:0]    _zz_sbuf_wdat_9_10;
  wire       [41:0]   _zz_sbuf_wdat_9_11;
  wire       [0:0]    _zz_sbuf_wdat_9_12;
  wire       [37:0]   _zz_sbuf_wdat_9_13;
  wire       [0:0]    _zz_sbuf_wdat_9_14;
  wire       [33:0]   _zz_sbuf_wdat_9_15;
  wire       [0:0]    _zz_sbuf_wdat_9_16;
  wire       [29:0]   _zz_sbuf_wdat_9_17;
  wire       [0:0]    _zz_sbuf_wdat_9_18;
  wire       [25:0]   _zz_sbuf_wdat_9_19;
  wire       [0:0]    _zz_sbuf_wdat_9_20;
  wire       [21:0]   _zz_sbuf_wdat_9_21;
  wire       [0:0]    _zz_sbuf_wdat_9_22;
  wire       [17:0]   _zz_sbuf_wdat_9_23;
  wire       [0:0]    _zz_sbuf_wdat_9_24;
  wire       [13:0]   _zz_sbuf_wdat_9_25;
  wire       [0:0]    _zz_sbuf_wdat_9_26;
  wire       [9:0]    _zz_sbuf_wdat_9_27;
  wire       [0:0]    _zz_sbuf_wdat_9_28;
  wire       [5:0]    _zz_sbuf_wdat_9_29;
  wire       [0:0]    _zz_sbuf_wdat_9_30;
  wire       [0:0]    _zz_sbuf_wdat_9_31;
  wire       [0:0]    _zz_sbuf_wdat_9_32;
  wire       [61:0]   _zz_sbuf_wdat_9_33;
  wire       [0:0]    _zz_sbuf_wdat_9_34;
  wire       [57:0]   _zz_sbuf_wdat_9_35;
  wire       [0:0]    _zz_sbuf_wdat_9_36;
  wire       [53:0]   _zz_sbuf_wdat_9_37;
  wire       [0:0]    _zz_sbuf_wdat_9_38;
  wire       [49:0]   _zz_sbuf_wdat_9_39;
  wire       [0:0]    _zz_sbuf_wdat_9_40;
  wire       [45:0]   _zz_sbuf_wdat_9_41;
  wire       [0:0]    _zz_sbuf_wdat_9_42;
  wire       [41:0]   _zz_sbuf_wdat_9_43;
  wire       [0:0]    _zz_sbuf_wdat_9_44;
  wire       [37:0]   _zz_sbuf_wdat_9_45;
  wire       [0:0]    _zz_sbuf_wdat_9_46;
  wire       [33:0]   _zz_sbuf_wdat_9_47;
  wire       [0:0]    _zz_sbuf_wdat_9_48;
  wire       [29:0]   _zz_sbuf_wdat_9_49;
  wire       [0:0]    _zz_sbuf_wdat_9_50;
  wire       [25:0]   _zz_sbuf_wdat_9_51;
  wire       [0:0]    _zz_sbuf_wdat_9_52;
  wire       [21:0]   _zz_sbuf_wdat_9_53;
  wire       [0:0]    _zz_sbuf_wdat_9_54;
  wire       [17:0]   _zz_sbuf_wdat_9_55;
  wire       [0:0]    _zz_sbuf_wdat_9_56;
  wire       [13:0]   _zz_sbuf_wdat_9_57;
  wire       [0:0]    _zz_sbuf_wdat_9_58;
  wire       [9:0]    _zz_sbuf_wdat_9_59;
  wire       [0:0]    _zz_sbuf_wdat_9_60;
  wire       [5:0]    _zz_sbuf_wdat_9_61;
  wire       [0:0]    _zz_sbuf_wdat_9_62;
  wire       [0:0]    _zz_sbuf_wdat_9_63;
  wire       [0:0]    _zz_sbuf_wdat_9_64;
  wire       [60:0]   _zz_sbuf_wdat_9_65;
  wire       [0:0]    _zz_sbuf_wdat_9_66;
  wire       [56:0]   _zz_sbuf_wdat_9_67;
  wire       [0:0]    _zz_sbuf_wdat_9_68;
  wire       [52:0]   _zz_sbuf_wdat_9_69;
  wire       [0:0]    _zz_sbuf_wdat_9_70;
  wire       [48:0]   _zz_sbuf_wdat_9_71;
  wire       [0:0]    _zz_sbuf_wdat_9_72;
  wire       [44:0]   _zz_sbuf_wdat_9_73;
  wire       [0:0]    _zz_sbuf_wdat_9_74;
  wire       [40:0]   _zz_sbuf_wdat_9_75;
  wire       [0:0]    _zz_sbuf_wdat_9_76;
  wire       [36:0]   _zz_sbuf_wdat_9_77;
  wire       [0:0]    _zz_sbuf_wdat_9_78;
  wire       [32:0]   _zz_sbuf_wdat_9_79;
  wire       [0:0]    _zz_sbuf_wdat_9_80;
  wire       [28:0]   _zz_sbuf_wdat_9_81;
  wire       [0:0]    _zz_sbuf_wdat_9_82;
  wire       [24:0]   _zz_sbuf_wdat_9_83;
  wire       [0:0]    _zz_sbuf_wdat_9_84;
  wire       [20:0]   _zz_sbuf_wdat_9_85;
  wire       [0:0]    _zz_sbuf_wdat_9_86;
  wire       [16:0]   _zz_sbuf_wdat_9_87;
  wire       [0:0]    _zz_sbuf_wdat_9_88;
  wire       [12:0]   _zz_sbuf_wdat_9_89;
  wire       [0:0]    _zz_sbuf_wdat_9_90;
  wire       [8:0]    _zz_sbuf_wdat_9_91;
  wire       [0:0]    _zz_sbuf_wdat_9_92;
  wire       [4:0]    _zz_sbuf_wdat_9_93;
  wire       [0:0]    _zz_sbuf_wdat_9_94;
  wire       [59:0]   _zz_sbuf_wdat_9_95;
  wire       [0:0]    _zz_sbuf_wdat_9_96;
  wire       [55:0]   _zz_sbuf_wdat_9_97;
  wire       [0:0]    _zz_sbuf_wdat_9_98;
  wire       [51:0]   _zz_sbuf_wdat_9_99;
  wire       [0:0]    _zz_sbuf_wdat_9_100;
  wire       [47:0]   _zz_sbuf_wdat_9_101;
  wire       [0:0]    _zz_sbuf_wdat_9_102;
  wire       [43:0]   _zz_sbuf_wdat_9_103;
  wire       [0:0]    _zz_sbuf_wdat_9_104;
  wire       [39:0]   _zz_sbuf_wdat_9_105;
  wire       [0:0]    _zz_sbuf_wdat_9_106;
  wire       [35:0]   _zz_sbuf_wdat_9_107;
  wire       [0:0]    _zz_sbuf_wdat_9_108;
  wire       [31:0]   _zz_sbuf_wdat_9_109;
  wire       [0:0]    _zz_sbuf_wdat_9_110;
  wire       [27:0]   _zz_sbuf_wdat_9_111;
  wire       [0:0]    _zz_sbuf_wdat_9_112;
  wire       [23:0]   _zz_sbuf_wdat_9_113;
  wire       [0:0]    _zz_sbuf_wdat_9_114;
  wire       [19:0]   _zz_sbuf_wdat_9_115;
  wire       [0:0]    _zz_sbuf_wdat_9_116;
  wire       [15:0]   _zz_sbuf_wdat_9_117;
  wire       [0:0]    _zz_sbuf_wdat_9_118;
  wire       [11:0]   _zz_sbuf_wdat_9_119;
  wire       [0:0]    _zz_sbuf_wdat_9_120;
  wire       [7:0]    _zz_sbuf_wdat_9_121;
  wire       [0:0]    _zz_sbuf_wdat_9_122;
  wire       [3:0]    _zz_sbuf_wdat_9_123;
  wire       [0:0]    _zz_sbuf_wdat_10;
  wire       [61:0]   _zz_sbuf_wdat_10_1;
  wire       [0:0]    _zz_sbuf_wdat_10_2;
  wire       [57:0]   _zz_sbuf_wdat_10_3;
  wire       [0:0]    _zz_sbuf_wdat_10_4;
  wire       [53:0]   _zz_sbuf_wdat_10_5;
  wire       [0:0]    _zz_sbuf_wdat_10_6;
  wire       [49:0]   _zz_sbuf_wdat_10_7;
  wire       [0:0]    _zz_sbuf_wdat_10_8;
  wire       [45:0]   _zz_sbuf_wdat_10_9;
  wire       [0:0]    _zz_sbuf_wdat_10_10;
  wire       [41:0]   _zz_sbuf_wdat_10_11;
  wire       [0:0]    _zz_sbuf_wdat_10_12;
  wire       [37:0]   _zz_sbuf_wdat_10_13;
  wire       [0:0]    _zz_sbuf_wdat_10_14;
  wire       [33:0]   _zz_sbuf_wdat_10_15;
  wire       [0:0]    _zz_sbuf_wdat_10_16;
  wire       [29:0]   _zz_sbuf_wdat_10_17;
  wire       [0:0]    _zz_sbuf_wdat_10_18;
  wire       [25:0]   _zz_sbuf_wdat_10_19;
  wire       [0:0]    _zz_sbuf_wdat_10_20;
  wire       [21:0]   _zz_sbuf_wdat_10_21;
  wire       [0:0]    _zz_sbuf_wdat_10_22;
  wire       [17:0]   _zz_sbuf_wdat_10_23;
  wire       [0:0]    _zz_sbuf_wdat_10_24;
  wire       [13:0]   _zz_sbuf_wdat_10_25;
  wire       [0:0]    _zz_sbuf_wdat_10_26;
  wire       [9:0]    _zz_sbuf_wdat_10_27;
  wire       [0:0]    _zz_sbuf_wdat_10_28;
  wire       [5:0]    _zz_sbuf_wdat_10_29;
  wire       [0:0]    _zz_sbuf_wdat_10_30;
  wire       [0:0]    _zz_sbuf_wdat_10_31;
  wire       [0:0]    _zz_sbuf_wdat_10_32;
  wire       [61:0]   _zz_sbuf_wdat_10_33;
  wire       [0:0]    _zz_sbuf_wdat_10_34;
  wire       [57:0]   _zz_sbuf_wdat_10_35;
  wire       [0:0]    _zz_sbuf_wdat_10_36;
  wire       [53:0]   _zz_sbuf_wdat_10_37;
  wire       [0:0]    _zz_sbuf_wdat_10_38;
  wire       [49:0]   _zz_sbuf_wdat_10_39;
  wire       [0:0]    _zz_sbuf_wdat_10_40;
  wire       [45:0]   _zz_sbuf_wdat_10_41;
  wire       [0:0]    _zz_sbuf_wdat_10_42;
  wire       [41:0]   _zz_sbuf_wdat_10_43;
  wire       [0:0]    _zz_sbuf_wdat_10_44;
  wire       [37:0]   _zz_sbuf_wdat_10_45;
  wire       [0:0]    _zz_sbuf_wdat_10_46;
  wire       [33:0]   _zz_sbuf_wdat_10_47;
  wire       [0:0]    _zz_sbuf_wdat_10_48;
  wire       [29:0]   _zz_sbuf_wdat_10_49;
  wire       [0:0]    _zz_sbuf_wdat_10_50;
  wire       [25:0]   _zz_sbuf_wdat_10_51;
  wire       [0:0]    _zz_sbuf_wdat_10_52;
  wire       [21:0]   _zz_sbuf_wdat_10_53;
  wire       [0:0]    _zz_sbuf_wdat_10_54;
  wire       [17:0]   _zz_sbuf_wdat_10_55;
  wire       [0:0]    _zz_sbuf_wdat_10_56;
  wire       [13:0]   _zz_sbuf_wdat_10_57;
  wire       [0:0]    _zz_sbuf_wdat_10_58;
  wire       [9:0]    _zz_sbuf_wdat_10_59;
  wire       [0:0]    _zz_sbuf_wdat_10_60;
  wire       [5:0]    _zz_sbuf_wdat_10_61;
  wire       [0:0]    _zz_sbuf_wdat_10_62;
  wire       [0:0]    _zz_sbuf_wdat_10_63;
  wire       [0:0]    _zz_sbuf_wdat_10_64;
  wire       [60:0]   _zz_sbuf_wdat_10_65;
  wire       [0:0]    _zz_sbuf_wdat_10_66;
  wire       [56:0]   _zz_sbuf_wdat_10_67;
  wire       [0:0]    _zz_sbuf_wdat_10_68;
  wire       [52:0]   _zz_sbuf_wdat_10_69;
  wire       [0:0]    _zz_sbuf_wdat_10_70;
  wire       [48:0]   _zz_sbuf_wdat_10_71;
  wire       [0:0]    _zz_sbuf_wdat_10_72;
  wire       [44:0]   _zz_sbuf_wdat_10_73;
  wire       [0:0]    _zz_sbuf_wdat_10_74;
  wire       [40:0]   _zz_sbuf_wdat_10_75;
  wire       [0:0]    _zz_sbuf_wdat_10_76;
  wire       [36:0]   _zz_sbuf_wdat_10_77;
  wire       [0:0]    _zz_sbuf_wdat_10_78;
  wire       [32:0]   _zz_sbuf_wdat_10_79;
  wire       [0:0]    _zz_sbuf_wdat_10_80;
  wire       [28:0]   _zz_sbuf_wdat_10_81;
  wire       [0:0]    _zz_sbuf_wdat_10_82;
  wire       [24:0]   _zz_sbuf_wdat_10_83;
  wire       [0:0]    _zz_sbuf_wdat_10_84;
  wire       [20:0]   _zz_sbuf_wdat_10_85;
  wire       [0:0]    _zz_sbuf_wdat_10_86;
  wire       [16:0]   _zz_sbuf_wdat_10_87;
  wire       [0:0]    _zz_sbuf_wdat_10_88;
  wire       [12:0]   _zz_sbuf_wdat_10_89;
  wire       [0:0]    _zz_sbuf_wdat_10_90;
  wire       [8:0]    _zz_sbuf_wdat_10_91;
  wire       [0:0]    _zz_sbuf_wdat_10_92;
  wire       [4:0]    _zz_sbuf_wdat_10_93;
  wire       [0:0]    _zz_sbuf_wdat_10_94;
  wire       [59:0]   _zz_sbuf_wdat_10_95;
  wire       [0:0]    _zz_sbuf_wdat_10_96;
  wire       [55:0]   _zz_sbuf_wdat_10_97;
  wire       [0:0]    _zz_sbuf_wdat_10_98;
  wire       [51:0]   _zz_sbuf_wdat_10_99;
  wire       [0:0]    _zz_sbuf_wdat_10_100;
  wire       [47:0]   _zz_sbuf_wdat_10_101;
  wire       [0:0]    _zz_sbuf_wdat_10_102;
  wire       [43:0]   _zz_sbuf_wdat_10_103;
  wire       [0:0]    _zz_sbuf_wdat_10_104;
  wire       [39:0]   _zz_sbuf_wdat_10_105;
  wire       [0:0]    _zz_sbuf_wdat_10_106;
  wire       [35:0]   _zz_sbuf_wdat_10_107;
  wire       [0:0]    _zz_sbuf_wdat_10_108;
  wire       [31:0]   _zz_sbuf_wdat_10_109;
  wire       [0:0]    _zz_sbuf_wdat_10_110;
  wire       [27:0]   _zz_sbuf_wdat_10_111;
  wire       [0:0]    _zz_sbuf_wdat_10_112;
  wire       [23:0]   _zz_sbuf_wdat_10_113;
  wire       [0:0]    _zz_sbuf_wdat_10_114;
  wire       [19:0]   _zz_sbuf_wdat_10_115;
  wire       [0:0]    _zz_sbuf_wdat_10_116;
  wire       [15:0]   _zz_sbuf_wdat_10_117;
  wire       [0:0]    _zz_sbuf_wdat_10_118;
  wire       [11:0]   _zz_sbuf_wdat_10_119;
  wire       [0:0]    _zz_sbuf_wdat_10_120;
  wire       [7:0]    _zz_sbuf_wdat_10_121;
  wire       [0:0]    _zz_sbuf_wdat_10_122;
  wire       [3:0]    _zz_sbuf_wdat_10_123;
  wire       [0:0]    _zz_sbuf_wdat_11;
  wire       [61:0]   _zz_sbuf_wdat_11_1;
  wire       [0:0]    _zz_sbuf_wdat_11_2;
  wire       [57:0]   _zz_sbuf_wdat_11_3;
  wire       [0:0]    _zz_sbuf_wdat_11_4;
  wire       [53:0]   _zz_sbuf_wdat_11_5;
  wire       [0:0]    _zz_sbuf_wdat_11_6;
  wire       [49:0]   _zz_sbuf_wdat_11_7;
  wire       [0:0]    _zz_sbuf_wdat_11_8;
  wire       [45:0]   _zz_sbuf_wdat_11_9;
  wire       [0:0]    _zz_sbuf_wdat_11_10;
  wire       [41:0]   _zz_sbuf_wdat_11_11;
  wire       [0:0]    _zz_sbuf_wdat_11_12;
  wire       [37:0]   _zz_sbuf_wdat_11_13;
  wire       [0:0]    _zz_sbuf_wdat_11_14;
  wire       [33:0]   _zz_sbuf_wdat_11_15;
  wire       [0:0]    _zz_sbuf_wdat_11_16;
  wire       [29:0]   _zz_sbuf_wdat_11_17;
  wire       [0:0]    _zz_sbuf_wdat_11_18;
  wire       [25:0]   _zz_sbuf_wdat_11_19;
  wire       [0:0]    _zz_sbuf_wdat_11_20;
  wire       [21:0]   _zz_sbuf_wdat_11_21;
  wire       [0:0]    _zz_sbuf_wdat_11_22;
  wire       [17:0]   _zz_sbuf_wdat_11_23;
  wire       [0:0]    _zz_sbuf_wdat_11_24;
  wire       [13:0]   _zz_sbuf_wdat_11_25;
  wire       [0:0]    _zz_sbuf_wdat_11_26;
  wire       [9:0]    _zz_sbuf_wdat_11_27;
  wire       [0:0]    _zz_sbuf_wdat_11_28;
  wire       [5:0]    _zz_sbuf_wdat_11_29;
  wire       [0:0]    _zz_sbuf_wdat_11_30;
  wire       [0:0]    _zz_sbuf_wdat_11_31;
  wire       [0:0]    _zz_sbuf_wdat_11_32;
  wire       [61:0]   _zz_sbuf_wdat_11_33;
  wire       [0:0]    _zz_sbuf_wdat_11_34;
  wire       [57:0]   _zz_sbuf_wdat_11_35;
  wire       [0:0]    _zz_sbuf_wdat_11_36;
  wire       [53:0]   _zz_sbuf_wdat_11_37;
  wire       [0:0]    _zz_sbuf_wdat_11_38;
  wire       [49:0]   _zz_sbuf_wdat_11_39;
  wire       [0:0]    _zz_sbuf_wdat_11_40;
  wire       [45:0]   _zz_sbuf_wdat_11_41;
  wire       [0:0]    _zz_sbuf_wdat_11_42;
  wire       [41:0]   _zz_sbuf_wdat_11_43;
  wire       [0:0]    _zz_sbuf_wdat_11_44;
  wire       [37:0]   _zz_sbuf_wdat_11_45;
  wire       [0:0]    _zz_sbuf_wdat_11_46;
  wire       [33:0]   _zz_sbuf_wdat_11_47;
  wire       [0:0]    _zz_sbuf_wdat_11_48;
  wire       [29:0]   _zz_sbuf_wdat_11_49;
  wire       [0:0]    _zz_sbuf_wdat_11_50;
  wire       [25:0]   _zz_sbuf_wdat_11_51;
  wire       [0:0]    _zz_sbuf_wdat_11_52;
  wire       [21:0]   _zz_sbuf_wdat_11_53;
  wire       [0:0]    _zz_sbuf_wdat_11_54;
  wire       [17:0]   _zz_sbuf_wdat_11_55;
  wire       [0:0]    _zz_sbuf_wdat_11_56;
  wire       [13:0]   _zz_sbuf_wdat_11_57;
  wire       [0:0]    _zz_sbuf_wdat_11_58;
  wire       [9:0]    _zz_sbuf_wdat_11_59;
  wire       [0:0]    _zz_sbuf_wdat_11_60;
  wire       [5:0]    _zz_sbuf_wdat_11_61;
  wire       [0:0]    _zz_sbuf_wdat_11_62;
  wire       [0:0]    _zz_sbuf_wdat_11_63;
  wire       [0:0]    _zz_sbuf_wdat_11_64;
  wire       [60:0]   _zz_sbuf_wdat_11_65;
  wire       [0:0]    _zz_sbuf_wdat_11_66;
  wire       [56:0]   _zz_sbuf_wdat_11_67;
  wire       [0:0]    _zz_sbuf_wdat_11_68;
  wire       [52:0]   _zz_sbuf_wdat_11_69;
  wire       [0:0]    _zz_sbuf_wdat_11_70;
  wire       [48:0]   _zz_sbuf_wdat_11_71;
  wire       [0:0]    _zz_sbuf_wdat_11_72;
  wire       [44:0]   _zz_sbuf_wdat_11_73;
  wire       [0:0]    _zz_sbuf_wdat_11_74;
  wire       [40:0]   _zz_sbuf_wdat_11_75;
  wire       [0:0]    _zz_sbuf_wdat_11_76;
  wire       [36:0]   _zz_sbuf_wdat_11_77;
  wire       [0:0]    _zz_sbuf_wdat_11_78;
  wire       [32:0]   _zz_sbuf_wdat_11_79;
  wire       [0:0]    _zz_sbuf_wdat_11_80;
  wire       [28:0]   _zz_sbuf_wdat_11_81;
  wire       [0:0]    _zz_sbuf_wdat_11_82;
  wire       [24:0]   _zz_sbuf_wdat_11_83;
  wire       [0:0]    _zz_sbuf_wdat_11_84;
  wire       [20:0]   _zz_sbuf_wdat_11_85;
  wire       [0:0]    _zz_sbuf_wdat_11_86;
  wire       [16:0]   _zz_sbuf_wdat_11_87;
  wire       [0:0]    _zz_sbuf_wdat_11_88;
  wire       [12:0]   _zz_sbuf_wdat_11_89;
  wire       [0:0]    _zz_sbuf_wdat_11_90;
  wire       [8:0]    _zz_sbuf_wdat_11_91;
  wire       [0:0]    _zz_sbuf_wdat_11_92;
  wire       [4:0]    _zz_sbuf_wdat_11_93;
  wire       [0:0]    _zz_sbuf_wdat_11_94;
  wire       [59:0]   _zz_sbuf_wdat_11_95;
  wire       [0:0]    _zz_sbuf_wdat_11_96;
  wire       [55:0]   _zz_sbuf_wdat_11_97;
  wire       [0:0]    _zz_sbuf_wdat_11_98;
  wire       [51:0]   _zz_sbuf_wdat_11_99;
  wire       [0:0]    _zz_sbuf_wdat_11_100;
  wire       [47:0]   _zz_sbuf_wdat_11_101;
  wire       [0:0]    _zz_sbuf_wdat_11_102;
  wire       [43:0]   _zz_sbuf_wdat_11_103;
  wire       [0:0]    _zz_sbuf_wdat_11_104;
  wire       [39:0]   _zz_sbuf_wdat_11_105;
  wire       [0:0]    _zz_sbuf_wdat_11_106;
  wire       [35:0]   _zz_sbuf_wdat_11_107;
  wire       [0:0]    _zz_sbuf_wdat_11_108;
  wire       [31:0]   _zz_sbuf_wdat_11_109;
  wire       [0:0]    _zz_sbuf_wdat_11_110;
  wire       [27:0]   _zz_sbuf_wdat_11_111;
  wire       [0:0]    _zz_sbuf_wdat_11_112;
  wire       [23:0]   _zz_sbuf_wdat_11_113;
  wire       [0:0]    _zz_sbuf_wdat_11_114;
  wire       [19:0]   _zz_sbuf_wdat_11_115;
  wire       [0:0]    _zz_sbuf_wdat_11_116;
  wire       [15:0]   _zz_sbuf_wdat_11_117;
  wire       [0:0]    _zz_sbuf_wdat_11_118;
  wire       [11:0]   _zz_sbuf_wdat_11_119;
  wire       [0:0]    _zz_sbuf_wdat_11_120;
  wire       [7:0]    _zz_sbuf_wdat_11_121;
  wire       [0:0]    _zz_sbuf_wdat_11_122;
  wire       [3:0]    _zz_sbuf_wdat_11_123;
  wire       [0:0]    _zz_sbuf_wdat_12;
  wire       [61:0]   _zz_sbuf_wdat_12_1;
  wire       [0:0]    _zz_sbuf_wdat_12_2;
  wire       [57:0]   _zz_sbuf_wdat_12_3;
  wire       [0:0]    _zz_sbuf_wdat_12_4;
  wire       [53:0]   _zz_sbuf_wdat_12_5;
  wire       [0:0]    _zz_sbuf_wdat_12_6;
  wire       [49:0]   _zz_sbuf_wdat_12_7;
  wire       [0:0]    _zz_sbuf_wdat_12_8;
  wire       [45:0]   _zz_sbuf_wdat_12_9;
  wire       [0:0]    _zz_sbuf_wdat_12_10;
  wire       [41:0]   _zz_sbuf_wdat_12_11;
  wire       [0:0]    _zz_sbuf_wdat_12_12;
  wire       [37:0]   _zz_sbuf_wdat_12_13;
  wire       [0:0]    _zz_sbuf_wdat_12_14;
  wire       [33:0]   _zz_sbuf_wdat_12_15;
  wire       [0:0]    _zz_sbuf_wdat_12_16;
  wire       [29:0]   _zz_sbuf_wdat_12_17;
  wire       [0:0]    _zz_sbuf_wdat_12_18;
  wire       [25:0]   _zz_sbuf_wdat_12_19;
  wire       [0:0]    _zz_sbuf_wdat_12_20;
  wire       [21:0]   _zz_sbuf_wdat_12_21;
  wire       [0:0]    _zz_sbuf_wdat_12_22;
  wire       [17:0]   _zz_sbuf_wdat_12_23;
  wire       [0:0]    _zz_sbuf_wdat_12_24;
  wire       [13:0]   _zz_sbuf_wdat_12_25;
  wire       [0:0]    _zz_sbuf_wdat_12_26;
  wire       [9:0]    _zz_sbuf_wdat_12_27;
  wire       [0:0]    _zz_sbuf_wdat_12_28;
  wire       [5:0]    _zz_sbuf_wdat_12_29;
  wire       [0:0]    _zz_sbuf_wdat_12_30;
  wire       [0:0]    _zz_sbuf_wdat_12_31;
  wire       [0:0]    _zz_sbuf_wdat_12_32;
  wire       [61:0]   _zz_sbuf_wdat_12_33;
  wire       [0:0]    _zz_sbuf_wdat_12_34;
  wire       [57:0]   _zz_sbuf_wdat_12_35;
  wire       [0:0]    _zz_sbuf_wdat_12_36;
  wire       [53:0]   _zz_sbuf_wdat_12_37;
  wire       [0:0]    _zz_sbuf_wdat_12_38;
  wire       [49:0]   _zz_sbuf_wdat_12_39;
  wire       [0:0]    _zz_sbuf_wdat_12_40;
  wire       [45:0]   _zz_sbuf_wdat_12_41;
  wire       [0:0]    _zz_sbuf_wdat_12_42;
  wire       [41:0]   _zz_sbuf_wdat_12_43;
  wire       [0:0]    _zz_sbuf_wdat_12_44;
  wire       [37:0]   _zz_sbuf_wdat_12_45;
  wire       [0:0]    _zz_sbuf_wdat_12_46;
  wire       [33:0]   _zz_sbuf_wdat_12_47;
  wire       [0:0]    _zz_sbuf_wdat_12_48;
  wire       [29:0]   _zz_sbuf_wdat_12_49;
  wire       [0:0]    _zz_sbuf_wdat_12_50;
  wire       [25:0]   _zz_sbuf_wdat_12_51;
  wire       [0:0]    _zz_sbuf_wdat_12_52;
  wire       [21:0]   _zz_sbuf_wdat_12_53;
  wire       [0:0]    _zz_sbuf_wdat_12_54;
  wire       [17:0]   _zz_sbuf_wdat_12_55;
  wire       [0:0]    _zz_sbuf_wdat_12_56;
  wire       [13:0]   _zz_sbuf_wdat_12_57;
  wire       [0:0]    _zz_sbuf_wdat_12_58;
  wire       [9:0]    _zz_sbuf_wdat_12_59;
  wire       [0:0]    _zz_sbuf_wdat_12_60;
  wire       [5:0]    _zz_sbuf_wdat_12_61;
  wire       [0:0]    _zz_sbuf_wdat_12_62;
  wire       [0:0]    _zz_sbuf_wdat_12_63;
  wire       [0:0]    _zz_sbuf_wdat_12_64;
  wire       [60:0]   _zz_sbuf_wdat_12_65;
  wire       [0:0]    _zz_sbuf_wdat_12_66;
  wire       [56:0]   _zz_sbuf_wdat_12_67;
  wire       [0:0]    _zz_sbuf_wdat_12_68;
  wire       [52:0]   _zz_sbuf_wdat_12_69;
  wire       [0:0]    _zz_sbuf_wdat_12_70;
  wire       [48:0]   _zz_sbuf_wdat_12_71;
  wire       [0:0]    _zz_sbuf_wdat_12_72;
  wire       [44:0]   _zz_sbuf_wdat_12_73;
  wire       [0:0]    _zz_sbuf_wdat_12_74;
  wire       [40:0]   _zz_sbuf_wdat_12_75;
  wire       [0:0]    _zz_sbuf_wdat_12_76;
  wire       [36:0]   _zz_sbuf_wdat_12_77;
  wire       [0:0]    _zz_sbuf_wdat_12_78;
  wire       [32:0]   _zz_sbuf_wdat_12_79;
  wire       [0:0]    _zz_sbuf_wdat_12_80;
  wire       [28:0]   _zz_sbuf_wdat_12_81;
  wire       [0:0]    _zz_sbuf_wdat_12_82;
  wire       [24:0]   _zz_sbuf_wdat_12_83;
  wire       [0:0]    _zz_sbuf_wdat_12_84;
  wire       [20:0]   _zz_sbuf_wdat_12_85;
  wire       [0:0]    _zz_sbuf_wdat_12_86;
  wire       [16:0]   _zz_sbuf_wdat_12_87;
  wire       [0:0]    _zz_sbuf_wdat_12_88;
  wire       [12:0]   _zz_sbuf_wdat_12_89;
  wire       [0:0]    _zz_sbuf_wdat_12_90;
  wire       [8:0]    _zz_sbuf_wdat_12_91;
  wire       [0:0]    _zz_sbuf_wdat_12_92;
  wire       [4:0]    _zz_sbuf_wdat_12_93;
  wire       [0:0]    _zz_sbuf_wdat_12_94;
  wire       [59:0]   _zz_sbuf_wdat_12_95;
  wire       [0:0]    _zz_sbuf_wdat_12_96;
  wire       [55:0]   _zz_sbuf_wdat_12_97;
  wire       [0:0]    _zz_sbuf_wdat_12_98;
  wire       [51:0]   _zz_sbuf_wdat_12_99;
  wire       [0:0]    _zz_sbuf_wdat_12_100;
  wire       [47:0]   _zz_sbuf_wdat_12_101;
  wire       [0:0]    _zz_sbuf_wdat_12_102;
  wire       [43:0]   _zz_sbuf_wdat_12_103;
  wire       [0:0]    _zz_sbuf_wdat_12_104;
  wire       [39:0]   _zz_sbuf_wdat_12_105;
  wire       [0:0]    _zz_sbuf_wdat_12_106;
  wire       [35:0]   _zz_sbuf_wdat_12_107;
  wire       [0:0]    _zz_sbuf_wdat_12_108;
  wire       [31:0]   _zz_sbuf_wdat_12_109;
  wire       [0:0]    _zz_sbuf_wdat_12_110;
  wire       [27:0]   _zz_sbuf_wdat_12_111;
  wire       [0:0]    _zz_sbuf_wdat_12_112;
  wire       [23:0]   _zz_sbuf_wdat_12_113;
  wire       [0:0]    _zz_sbuf_wdat_12_114;
  wire       [19:0]   _zz_sbuf_wdat_12_115;
  wire       [0:0]    _zz_sbuf_wdat_12_116;
  wire       [15:0]   _zz_sbuf_wdat_12_117;
  wire       [0:0]    _zz_sbuf_wdat_12_118;
  wire       [11:0]   _zz_sbuf_wdat_12_119;
  wire       [0:0]    _zz_sbuf_wdat_12_120;
  wire       [7:0]    _zz_sbuf_wdat_12_121;
  wire       [0:0]    _zz_sbuf_wdat_12_122;
  wire       [3:0]    _zz_sbuf_wdat_12_123;
  wire       [0:0]    _zz_sbuf_wdat_13;
  wire       [61:0]   _zz_sbuf_wdat_13_1;
  wire       [0:0]    _zz_sbuf_wdat_13_2;
  wire       [57:0]   _zz_sbuf_wdat_13_3;
  wire       [0:0]    _zz_sbuf_wdat_13_4;
  wire       [53:0]   _zz_sbuf_wdat_13_5;
  wire       [0:0]    _zz_sbuf_wdat_13_6;
  wire       [49:0]   _zz_sbuf_wdat_13_7;
  wire       [0:0]    _zz_sbuf_wdat_13_8;
  wire       [45:0]   _zz_sbuf_wdat_13_9;
  wire       [0:0]    _zz_sbuf_wdat_13_10;
  wire       [41:0]   _zz_sbuf_wdat_13_11;
  wire       [0:0]    _zz_sbuf_wdat_13_12;
  wire       [37:0]   _zz_sbuf_wdat_13_13;
  wire       [0:0]    _zz_sbuf_wdat_13_14;
  wire       [33:0]   _zz_sbuf_wdat_13_15;
  wire       [0:0]    _zz_sbuf_wdat_13_16;
  wire       [29:0]   _zz_sbuf_wdat_13_17;
  wire       [0:0]    _zz_sbuf_wdat_13_18;
  wire       [25:0]   _zz_sbuf_wdat_13_19;
  wire       [0:0]    _zz_sbuf_wdat_13_20;
  wire       [21:0]   _zz_sbuf_wdat_13_21;
  wire       [0:0]    _zz_sbuf_wdat_13_22;
  wire       [17:0]   _zz_sbuf_wdat_13_23;
  wire       [0:0]    _zz_sbuf_wdat_13_24;
  wire       [13:0]   _zz_sbuf_wdat_13_25;
  wire       [0:0]    _zz_sbuf_wdat_13_26;
  wire       [9:0]    _zz_sbuf_wdat_13_27;
  wire       [0:0]    _zz_sbuf_wdat_13_28;
  wire       [5:0]    _zz_sbuf_wdat_13_29;
  wire       [0:0]    _zz_sbuf_wdat_13_30;
  wire       [0:0]    _zz_sbuf_wdat_13_31;
  wire       [0:0]    _zz_sbuf_wdat_13_32;
  wire       [61:0]   _zz_sbuf_wdat_13_33;
  wire       [0:0]    _zz_sbuf_wdat_13_34;
  wire       [57:0]   _zz_sbuf_wdat_13_35;
  wire       [0:0]    _zz_sbuf_wdat_13_36;
  wire       [53:0]   _zz_sbuf_wdat_13_37;
  wire       [0:0]    _zz_sbuf_wdat_13_38;
  wire       [49:0]   _zz_sbuf_wdat_13_39;
  wire       [0:0]    _zz_sbuf_wdat_13_40;
  wire       [45:0]   _zz_sbuf_wdat_13_41;
  wire       [0:0]    _zz_sbuf_wdat_13_42;
  wire       [41:0]   _zz_sbuf_wdat_13_43;
  wire       [0:0]    _zz_sbuf_wdat_13_44;
  wire       [37:0]   _zz_sbuf_wdat_13_45;
  wire       [0:0]    _zz_sbuf_wdat_13_46;
  wire       [33:0]   _zz_sbuf_wdat_13_47;
  wire       [0:0]    _zz_sbuf_wdat_13_48;
  wire       [29:0]   _zz_sbuf_wdat_13_49;
  wire       [0:0]    _zz_sbuf_wdat_13_50;
  wire       [25:0]   _zz_sbuf_wdat_13_51;
  wire       [0:0]    _zz_sbuf_wdat_13_52;
  wire       [21:0]   _zz_sbuf_wdat_13_53;
  wire       [0:0]    _zz_sbuf_wdat_13_54;
  wire       [17:0]   _zz_sbuf_wdat_13_55;
  wire       [0:0]    _zz_sbuf_wdat_13_56;
  wire       [13:0]   _zz_sbuf_wdat_13_57;
  wire       [0:0]    _zz_sbuf_wdat_13_58;
  wire       [9:0]    _zz_sbuf_wdat_13_59;
  wire       [0:0]    _zz_sbuf_wdat_13_60;
  wire       [5:0]    _zz_sbuf_wdat_13_61;
  wire       [0:0]    _zz_sbuf_wdat_13_62;
  wire       [0:0]    _zz_sbuf_wdat_13_63;
  wire       [0:0]    _zz_sbuf_wdat_13_64;
  wire       [60:0]   _zz_sbuf_wdat_13_65;
  wire       [0:0]    _zz_sbuf_wdat_13_66;
  wire       [56:0]   _zz_sbuf_wdat_13_67;
  wire       [0:0]    _zz_sbuf_wdat_13_68;
  wire       [52:0]   _zz_sbuf_wdat_13_69;
  wire       [0:0]    _zz_sbuf_wdat_13_70;
  wire       [48:0]   _zz_sbuf_wdat_13_71;
  wire       [0:0]    _zz_sbuf_wdat_13_72;
  wire       [44:0]   _zz_sbuf_wdat_13_73;
  wire       [0:0]    _zz_sbuf_wdat_13_74;
  wire       [40:0]   _zz_sbuf_wdat_13_75;
  wire       [0:0]    _zz_sbuf_wdat_13_76;
  wire       [36:0]   _zz_sbuf_wdat_13_77;
  wire       [0:0]    _zz_sbuf_wdat_13_78;
  wire       [32:0]   _zz_sbuf_wdat_13_79;
  wire       [0:0]    _zz_sbuf_wdat_13_80;
  wire       [28:0]   _zz_sbuf_wdat_13_81;
  wire       [0:0]    _zz_sbuf_wdat_13_82;
  wire       [24:0]   _zz_sbuf_wdat_13_83;
  wire       [0:0]    _zz_sbuf_wdat_13_84;
  wire       [20:0]   _zz_sbuf_wdat_13_85;
  wire       [0:0]    _zz_sbuf_wdat_13_86;
  wire       [16:0]   _zz_sbuf_wdat_13_87;
  wire       [0:0]    _zz_sbuf_wdat_13_88;
  wire       [12:0]   _zz_sbuf_wdat_13_89;
  wire       [0:0]    _zz_sbuf_wdat_13_90;
  wire       [8:0]    _zz_sbuf_wdat_13_91;
  wire       [0:0]    _zz_sbuf_wdat_13_92;
  wire       [4:0]    _zz_sbuf_wdat_13_93;
  wire       [0:0]    _zz_sbuf_wdat_13_94;
  wire       [59:0]   _zz_sbuf_wdat_13_95;
  wire       [0:0]    _zz_sbuf_wdat_13_96;
  wire       [55:0]   _zz_sbuf_wdat_13_97;
  wire       [0:0]    _zz_sbuf_wdat_13_98;
  wire       [51:0]   _zz_sbuf_wdat_13_99;
  wire       [0:0]    _zz_sbuf_wdat_13_100;
  wire       [47:0]   _zz_sbuf_wdat_13_101;
  wire       [0:0]    _zz_sbuf_wdat_13_102;
  wire       [43:0]   _zz_sbuf_wdat_13_103;
  wire       [0:0]    _zz_sbuf_wdat_13_104;
  wire       [39:0]   _zz_sbuf_wdat_13_105;
  wire       [0:0]    _zz_sbuf_wdat_13_106;
  wire       [35:0]   _zz_sbuf_wdat_13_107;
  wire       [0:0]    _zz_sbuf_wdat_13_108;
  wire       [31:0]   _zz_sbuf_wdat_13_109;
  wire       [0:0]    _zz_sbuf_wdat_13_110;
  wire       [27:0]   _zz_sbuf_wdat_13_111;
  wire       [0:0]    _zz_sbuf_wdat_13_112;
  wire       [23:0]   _zz_sbuf_wdat_13_113;
  wire       [0:0]    _zz_sbuf_wdat_13_114;
  wire       [19:0]   _zz_sbuf_wdat_13_115;
  wire       [0:0]    _zz_sbuf_wdat_13_116;
  wire       [15:0]   _zz_sbuf_wdat_13_117;
  wire       [0:0]    _zz_sbuf_wdat_13_118;
  wire       [11:0]   _zz_sbuf_wdat_13_119;
  wire       [0:0]    _zz_sbuf_wdat_13_120;
  wire       [7:0]    _zz_sbuf_wdat_13_121;
  wire       [0:0]    _zz_sbuf_wdat_13_122;
  wire       [3:0]    _zz_sbuf_wdat_13_123;
  wire       [0:0]    _zz_sbuf_wdat_14;
  wire       [61:0]   _zz_sbuf_wdat_14_1;
  wire       [0:0]    _zz_sbuf_wdat_14_2;
  wire       [57:0]   _zz_sbuf_wdat_14_3;
  wire       [0:0]    _zz_sbuf_wdat_14_4;
  wire       [53:0]   _zz_sbuf_wdat_14_5;
  wire       [0:0]    _zz_sbuf_wdat_14_6;
  wire       [49:0]   _zz_sbuf_wdat_14_7;
  wire       [0:0]    _zz_sbuf_wdat_14_8;
  wire       [45:0]   _zz_sbuf_wdat_14_9;
  wire       [0:0]    _zz_sbuf_wdat_14_10;
  wire       [41:0]   _zz_sbuf_wdat_14_11;
  wire       [0:0]    _zz_sbuf_wdat_14_12;
  wire       [37:0]   _zz_sbuf_wdat_14_13;
  wire       [0:0]    _zz_sbuf_wdat_14_14;
  wire       [33:0]   _zz_sbuf_wdat_14_15;
  wire       [0:0]    _zz_sbuf_wdat_14_16;
  wire       [29:0]   _zz_sbuf_wdat_14_17;
  wire       [0:0]    _zz_sbuf_wdat_14_18;
  wire       [25:0]   _zz_sbuf_wdat_14_19;
  wire       [0:0]    _zz_sbuf_wdat_14_20;
  wire       [21:0]   _zz_sbuf_wdat_14_21;
  wire       [0:0]    _zz_sbuf_wdat_14_22;
  wire       [17:0]   _zz_sbuf_wdat_14_23;
  wire       [0:0]    _zz_sbuf_wdat_14_24;
  wire       [13:0]   _zz_sbuf_wdat_14_25;
  wire       [0:0]    _zz_sbuf_wdat_14_26;
  wire       [9:0]    _zz_sbuf_wdat_14_27;
  wire       [0:0]    _zz_sbuf_wdat_14_28;
  wire       [5:0]    _zz_sbuf_wdat_14_29;
  wire       [0:0]    _zz_sbuf_wdat_14_30;
  wire       [0:0]    _zz_sbuf_wdat_14_31;
  wire       [0:0]    _zz_sbuf_wdat_14_32;
  wire       [61:0]   _zz_sbuf_wdat_14_33;
  wire       [0:0]    _zz_sbuf_wdat_14_34;
  wire       [57:0]   _zz_sbuf_wdat_14_35;
  wire       [0:0]    _zz_sbuf_wdat_14_36;
  wire       [53:0]   _zz_sbuf_wdat_14_37;
  wire       [0:0]    _zz_sbuf_wdat_14_38;
  wire       [49:0]   _zz_sbuf_wdat_14_39;
  wire       [0:0]    _zz_sbuf_wdat_14_40;
  wire       [45:0]   _zz_sbuf_wdat_14_41;
  wire       [0:0]    _zz_sbuf_wdat_14_42;
  wire       [41:0]   _zz_sbuf_wdat_14_43;
  wire       [0:0]    _zz_sbuf_wdat_14_44;
  wire       [37:0]   _zz_sbuf_wdat_14_45;
  wire       [0:0]    _zz_sbuf_wdat_14_46;
  wire       [33:0]   _zz_sbuf_wdat_14_47;
  wire       [0:0]    _zz_sbuf_wdat_14_48;
  wire       [29:0]   _zz_sbuf_wdat_14_49;
  wire       [0:0]    _zz_sbuf_wdat_14_50;
  wire       [25:0]   _zz_sbuf_wdat_14_51;
  wire       [0:0]    _zz_sbuf_wdat_14_52;
  wire       [21:0]   _zz_sbuf_wdat_14_53;
  wire       [0:0]    _zz_sbuf_wdat_14_54;
  wire       [17:0]   _zz_sbuf_wdat_14_55;
  wire       [0:0]    _zz_sbuf_wdat_14_56;
  wire       [13:0]   _zz_sbuf_wdat_14_57;
  wire       [0:0]    _zz_sbuf_wdat_14_58;
  wire       [9:0]    _zz_sbuf_wdat_14_59;
  wire       [0:0]    _zz_sbuf_wdat_14_60;
  wire       [5:0]    _zz_sbuf_wdat_14_61;
  wire       [0:0]    _zz_sbuf_wdat_14_62;
  wire       [0:0]    _zz_sbuf_wdat_14_63;
  wire       [0:0]    _zz_sbuf_wdat_14_64;
  wire       [60:0]   _zz_sbuf_wdat_14_65;
  wire       [0:0]    _zz_sbuf_wdat_14_66;
  wire       [56:0]   _zz_sbuf_wdat_14_67;
  wire       [0:0]    _zz_sbuf_wdat_14_68;
  wire       [52:0]   _zz_sbuf_wdat_14_69;
  wire       [0:0]    _zz_sbuf_wdat_14_70;
  wire       [48:0]   _zz_sbuf_wdat_14_71;
  wire       [0:0]    _zz_sbuf_wdat_14_72;
  wire       [44:0]   _zz_sbuf_wdat_14_73;
  wire       [0:0]    _zz_sbuf_wdat_14_74;
  wire       [40:0]   _zz_sbuf_wdat_14_75;
  wire       [0:0]    _zz_sbuf_wdat_14_76;
  wire       [36:0]   _zz_sbuf_wdat_14_77;
  wire       [0:0]    _zz_sbuf_wdat_14_78;
  wire       [32:0]   _zz_sbuf_wdat_14_79;
  wire       [0:0]    _zz_sbuf_wdat_14_80;
  wire       [28:0]   _zz_sbuf_wdat_14_81;
  wire       [0:0]    _zz_sbuf_wdat_14_82;
  wire       [24:0]   _zz_sbuf_wdat_14_83;
  wire       [0:0]    _zz_sbuf_wdat_14_84;
  wire       [20:0]   _zz_sbuf_wdat_14_85;
  wire       [0:0]    _zz_sbuf_wdat_14_86;
  wire       [16:0]   _zz_sbuf_wdat_14_87;
  wire       [0:0]    _zz_sbuf_wdat_14_88;
  wire       [12:0]   _zz_sbuf_wdat_14_89;
  wire       [0:0]    _zz_sbuf_wdat_14_90;
  wire       [8:0]    _zz_sbuf_wdat_14_91;
  wire       [0:0]    _zz_sbuf_wdat_14_92;
  wire       [4:0]    _zz_sbuf_wdat_14_93;
  wire       [0:0]    _zz_sbuf_wdat_14_94;
  wire       [59:0]   _zz_sbuf_wdat_14_95;
  wire       [0:0]    _zz_sbuf_wdat_14_96;
  wire       [55:0]   _zz_sbuf_wdat_14_97;
  wire       [0:0]    _zz_sbuf_wdat_14_98;
  wire       [51:0]   _zz_sbuf_wdat_14_99;
  wire       [0:0]    _zz_sbuf_wdat_14_100;
  wire       [47:0]   _zz_sbuf_wdat_14_101;
  wire       [0:0]    _zz_sbuf_wdat_14_102;
  wire       [43:0]   _zz_sbuf_wdat_14_103;
  wire       [0:0]    _zz_sbuf_wdat_14_104;
  wire       [39:0]   _zz_sbuf_wdat_14_105;
  wire       [0:0]    _zz_sbuf_wdat_14_106;
  wire       [35:0]   _zz_sbuf_wdat_14_107;
  wire       [0:0]    _zz_sbuf_wdat_14_108;
  wire       [31:0]   _zz_sbuf_wdat_14_109;
  wire       [0:0]    _zz_sbuf_wdat_14_110;
  wire       [27:0]   _zz_sbuf_wdat_14_111;
  wire       [0:0]    _zz_sbuf_wdat_14_112;
  wire       [23:0]   _zz_sbuf_wdat_14_113;
  wire       [0:0]    _zz_sbuf_wdat_14_114;
  wire       [19:0]   _zz_sbuf_wdat_14_115;
  wire       [0:0]    _zz_sbuf_wdat_14_116;
  wire       [15:0]   _zz_sbuf_wdat_14_117;
  wire       [0:0]    _zz_sbuf_wdat_14_118;
  wire       [11:0]   _zz_sbuf_wdat_14_119;
  wire       [0:0]    _zz_sbuf_wdat_14_120;
  wire       [7:0]    _zz_sbuf_wdat_14_121;
  wire       [0:0]    _zz_sbuf_wdat_14_122;
  wire       [3:0]    _zz_sbuf_wdat_14_123;
  wire       [0:0]    _zz_sbuf_wdat_15;
  wire       [61:0]   _zz_sbuf_wdat_15_1;
  wire       [0:0]    _zz_sbuf_wdat_15_2;
  wire       [57:0]   _zz_sbuf_wdat_15_3;
  wire       [0:0]    _zz_sbuf_wdat_15_4;
  wire       [53:0]   _zz_sbuf_wdat_15_5;
  wire       [0:0]    _zz_sbuf_wdat_15_6;
  wire       [49:0]   _zz_sbuf_wdat_15_7;
  wire       [0:0]    _zz_sbuf_wdat_15_8;
  wire       [45:0]   _zz_sbuf_wdat_15_9;
  wire       [0:0]    _zz_sbuf_wdat_15_10;
  wire       [41:0]   _zz_sbuf_wdat_15_11;
  wire       [0:0]    _zz_sbuf_wdat_15_12;
  wire       [37:0]   _zz_sbuf_wdat_15_13;
  wire       [0:0]    _zz_sbuf_wdat_15_14;
  wire       [33:0]   _zz_sbuf_wdat_15_15;
  wire       [0:0]    _zz_sbuf_wdat_15_16;
  wire       [29:0]   _zz_sbuf_wdat_15_17;
  wire       [0:0]    _zz_sbuf_wdat_15_18;
  wire       [25:0]   _zz_sbuf_wdat_15_19;
  wire       [0:0]    _zz_sbuf_wdat_15_20;
  wire       [21:0]   _zz_sbuf_wdat_15_21;
  wire       [0:0]    _zz_sbuf_wdat_15_22;
  wire       [17:0]   _zz_sbuf_wdat_15_23;
  wire       [0:0]    _zz_sbuf_wdat_15_24;
  wire       [13:0]   _zz_sbuf_wdat_15_25;
  wire       [0:0]    _zz_sbuf_wdat_15_26;
  wire       [9:0]    _zz_sbuf_wdat_15_27;
  wire       [0:0]    _zz_sbuf_wdat_15_28;
  wire       [5:0]    _zz_sbuf_wdat_15_29;
  wire       [0:0]    _zz_sbuf_wdat_15_30;
  wire       [0:0]    _zz_sbuf_wdat_15_31;
  wire       [0:0]    _zz_sbuf_wdat_15_32;
  wire       [61:0]   _zz_sbuf_wdat_15_33;
  wire       [0:0]    _zz_sbuf_wdat_15_34;
  wire       [57:0]   _zz_sbuf_wdat_15_35;
  wire       [0:0]    _zz_sbuf_wdat_15_36;
  wire       [53:0]   _zz_sbuf_wdat_15_37;
  wire       [0:0]    _zz_sbuf_wdat_15_38;
  wire       [49:0]   _zz_sbuf_wdat_15_39;
  wire       [0:0]    _zz_sbuf_wdat_15_40;
  wire       [45:0]   _zz_sbuf_wdat_15_41;
  wire       [0:0]    _zz_sbuf_wdat_15_42;
  wire       [41:0]   _zz_sbuf_wdat_15_43;
  wire       [0:0]    _zz_sbuf_wdat_15_44;
  wire       [37:0]   _zz_sbuf_wdat_15_45;
  wire       [0:0]    _zz_sbuf_wdat_15_46;
  wire       [33:0]   _zz_sbuf_wdat_15_47;
  wire       [0:0]    _zz_sbuf_wdat_15_48;
  wire       [29:0]   _zz_sbuf_wdat_15_49;
  wire       [0:0]    _zz_sbuf_wdat_15_50;
  wire       [25:0]   _zz_sbuf_wdat_15_51;
  wire       [0:0]    _zz_sbuf_wdat_15_52;
  wire       [21:0]   _zz_sbuf_wdat_15_53;
  wire       [0:0]    _zz_sbuf_wdat_15_54;
  wire       [17:0]   _zz_sbuf_wdat_15_55;
  wire       [0:0]    _zz_sbuf_wdat_15_56;
  wire       [13:0]   _zz_sbuf_wdat_15_57;
  wire       [0:0]    _zz_sbuf_wdat_15_58;
  wire       [9:0]    _zz_sbuf_wdat_15_59;
  wire       [0:0]    _zz_sbuf_wdat_15_60;
  wire       [5:0]    _zz_sbuf_wdat_15_61;
  wire       [0:0]    _zz_sbuf_wdat_15_62;
  wire       [0:0]    _zz_sbuf_wdat_15_63;
  wire       [0:0]    _zz_sbuf_wdat_15_64;
  wire       [60:0]   _zz_sbuf_wdat_15_65;
  wire       [0:0]    _zz_sbuf_wdat_15_66;
  wire       [56:0]   _zz_sbuf_wdat_15_67;
  wire       [0:0]    _zz_sbuf_wdat_15_68;
  wire       [52:0]   _zz_sbuf_wdat_15_69;
  wire       [0:0]    _zz_sbuf_wdat_15_70;
  wire       [48:0]   _zz_sbuf_wdat_15_71;
  wire       [0:0]    _zz_sbuf_wdat_15_72;
  wire       [44:0]   _zz_sbuf_wdat_15_73;
  wire       [0:0]    _zz_sbuf_wdat_15_74;
  wire       [40:0]   _zz_sbuf_wdat_15_75;
  wire       [0:0]    _zz_sbuf_wdat_15_76;
  wire       [36:0]   _zz_sbuf_wdat_15_77;
  wire       [0:0]    _zz_sbuf_wdat_15_78;
  wire       [32:0]   _zz_sbuf_wdat_15_79;
  wire       [0:0]    _zz_sbuf_wdat_15_80;
  wire       [28:0]   _zz_sbuf_wdat_15_81;
  wire       [0:0]    _zz_sbuf_wdat_15_82;
  wire       [24:0]   _zz_sbuf_wdat_15_83;
  wire       [0:0]    _zz_sbuf_wdat_15_84;
  wire       [20:0]   _zz_sbuf_wdat_15_85;
  wire       [0:0]    _zz_sbuf_wdat_15_86;
  wire       [16:0]   _zz_sbuf_wdat_15_87;
  wire       [0:0]    _zz_sbuf_wdat_15_88;
  wire       [12:0]   _zz_sbuf_wdat_15_89;
  wire       [0:0]    _zz_sbuf_wdat_15_90;
  wire       [8:0]    _zz_sbuf_wdat_15_91;
  wire       [0:0]    _zz_sbuf_wdat_15_92;
  wire       [4:0]    _zz_sbuf_wdat_15_93;
  wire       [0:0]    _zz_sbuf_wdat_15_94;
  wire       [59:0]   _zz_sbuf_wdat_15_95;
  wire       [0:0]    _zz_sbuf_wdat_15_96;
  wire       [55:0]   _zz_sbuf_wdat_15_97;
  wire       [0:0]    _zz_sbuf_wdat_15_98;
  wire       [51:0]   _zz_sbuf_wdat_15_99;
  wire       [0:0]    _zz_sbuf_wdat_15_100;
  wire       [47:0]   _zz_sbuf_wdat_15_101;
  wire       [0:0]    _zz_sbuf_wdat_15_102;
  wire       [43:0]   _zz_sbuf_wdat_15_103;
  wire       [0:0]    _zz_sbuf_wdat_15_104;
  wire       [39:0]   _zz_sbuf_wdat_15_105;
  wire       [0:0]    _zz_sbuf_wdat_15_106;
  wire       [35:0]   _zz_sbuf_wdat_15_107;
  wire       [0:0]    _zz_sbuf_wdat_15_108;
  wire       [31:0]   _zz_sbuf_wdat_15_109;
  wire       [0:0]    _zz_sbuf_wdat_15_110;
  wire       [27:0]   _zz_sbuf_wdat_15_111;
  wire       [0:0]    _zz_sbuf_wdat_15_112;
  wire       [23:0]   _zz_sbuf_wdat_15_113;
  wire       [0:0]    _zz_sbuf_wdat_15_114;
  wire       [19:0]   _zz_sbuf_wdat_15_115;
  wire       [0:0]    _zz_sbuf_wdat_15_116;
  wire       [15:0]   _zz_sbuf_wdat_15_117;
  wire       [0:0]    _zz_sbuf_wdat_15_118;
  wire       [11:0]   _zz_sbuf_wdat_15_119;
  wire       [0:0]    _zz_sbuf_wdat_15_120;
  wire       [7:0]    _zz_sbuf_wdat_15_121;
  wire       [0:0]    _zz_sbuf_wdat_15_122;
  wire       [3:0]    _zz_sbuf_wdat_15_123;
  wire       [0:0]    _zz_sbuf_ra_0;
  wire       [2:0]    _zz_sbuf_ra_0_1;
  wire       [3:0]    _zz_sbuf_ra_0_2;
  wire       [0:0]    _zz_sbuf_ra_0_3;
  wire       [2:0]    _zz_sbuf_ra_0_4;
  wire       [3:0]    _zz_sbuf_ra_0_5;
  wire       [0:0]    _zz_sbuf_ra_0_6;
  wire       [1:0]    _zz_sbuf_ra_0_7;
  wire       [0:0]    _zz_sbuf_ra_0_8;
  wire       [0:0]    _zz_sbuf_ra_0_9;
  wire       [0:0]    _zz_sbuf_ra_1;
  wire       [2:0]    _zz_sbuf_ra_1_1;
  wire       [3:0]    _zz_sbuf_ra_1_2;
  wire       [0:0]    _zz_sbuf_ra_1_3;
  wire       [2:0]    _zz_sbuf_ra_1_4;
  wire       [3:0]    _zz_sbuf_ra_1_5;
  wire       [0:0]    _zz_sbuf_ra_1_6;
  wire       [1:0]    _zz_sbuf_ra_1_7;
  wire       [0:0]    _zz_sbuf_ra_1_8;
  wire       [0:0]    _zz_sbuf_ra_1_9;
  wire       [0:0]    _zz_sbuf_ra_2;
  wire       [2:0]    _zz_sbuf_ra_2_1;
  wire       [3:0]    _zz_sbuf_ra_2_2;
  wire       [0:0]    _zz_sbuf_ra_2_3;
  wire       [2:0]    _zz_sbuf_ra_2_4;
  wire       [3:0]    _zz_sbuf_ra_2_5;
  wire       [0:0]    _zz_sbuf_ra_2_6;
  wire       [1:0]    _zz_sbuf_ra_2_7;
  wire       [0:0]    _zz_sbuf_ra_2_8;
  wire       [0:0]    _zz_sbuf_ra_2_9;
  wire       [0:0]    _zz_sbuf_ra_3;
  wire       [2:0]    _zz_sbuf_ra_3_1;
  wire       [3:0]    _zz_sbuf_ra_3_2;
  wire       [0:0]    _zz_sbuf_ra_3_3;
  wire       [2:0]    _zz_sbuf_ra_3_4;
  wire       [3:0]    _zz_sbuf_ra_3_5;
  wire       [0:0]    _zz_sbuf_ra_3_6;
  wire       [1:0]    _zz_sbuf_ra_3_7;
  wire       [0:0]    _zz_sbuf_ra_3_8;
  wire       [0:0]    _zz_sbuf_ra_3_9;
  wire       [0:0]    _zz_sbuf_ra_4;
  wire       [2:0]    _zz_sbuf_ra_4_1;
  wire       [3:0]    _zz_sbuf_ra_4_2;
  wire       [0:0]    _zz_sbuf_ra_4_3;
  wire       [2:0]    _zz_sbuf_ra_4_4;
  wire       [3:0]    _zz_sbuf_ra_4_5;
  wire       [0:0]    _zz_sbuf_ra_4_6;
  wire       [1:0]    _zz_sbuf_ra_4_7;
  wire       [0:0]    _zz_sbuf_ra_4_8;
  wire       [0:0]    _zz_sbuf_ra_4_9;
  wire       [0:0]    _zz_sbuf_ra_5;
  wire       [2:0]    _zz_sbuf_ra_5_1;
  wire       [3:0]    _zz_sbuf_ra_5_2;
  wire       [0:0]    _zz_sbuf_ra_5_3;
  wire       [2:0]    _zz_sbuf_ra_5_4;
  wire       [3:0]    _zz_sbuf_ra_5_5;
  wire       [0:0]    _zz_sbuf_ra_5_6;
  wire       [1:0]    _zz_sbuf_ra_5_7;
  wire       [0:0]    _zz_sbuf_ra_5_8;
  wire       [0:0]    _zz_sbuf_ra_5_9;
  wire       [0:0]    _zz_sbuf_ra_6;
  wire       [2:0]    _zz_sbuf_ra_6_1;
  wire       [3:0]    _zz_sbuf_ra_6_2;
  wire       [0:0]    _zz_sbuf_ra_6_3;
  wire       [2:0]    _zz_sbuf_ra_6_4;
  wire       [3:0]    _zz_sbuf_ra_6_5;
  wire       [0:0]    _zz_sbuf_ra_6_6;
  wire       [1:0]    _zz_sbuf_ra_6_7;
  wire       [0:0]    _zz_sbuf_ra_6_8;
  wire       [0:0]    _zz_sbuf_ra_6_9;
  wire       [0:0]    _zz_sbuf_ra_7;
  wire       [2:0]    _zz_sbuf_ra_7_1;
  wire       [3:0]    _zz_sbuf_ra_7_2;
  wire       [0:0]    _zz_sbuf_ra_7_3;
  wire       [2:0]    _zz_sbuf_ra_7_4;
  wire       [3:0]    _zz_sbuf_ra_7_5;
  wire       [0:0]    _zz_sbuf_ra_7_6;
  wire       [1:0]    _zz_sbuf_ra_7_7;
  wire       [0:0]    _zz_sbuf_ra_7_8;
  wire       [0:0]    _zz_sbuf_ra_7_9;
  wire       [0:0]    _zz_sbuf_ra_8;
  wire       [2:0]    _zz_sbuf_ra_8_1;
  wire       [3:0]    _zz_sbuf_ra_8_2;
  wire       [0:0]    _zz_sbuf_ra_8_3;
  wire       [2:0]    _zz_sbuf_ra_8_4;
  wire       [3:0]    _zz_sbuf_ra_8_5;
  wire       [0:0]    _zz_sbuf_ra_8_6;
  wire       [1:0]    _zz_sbuf_ra_8_7;
  wire       [0:0]    _zz_sbuf_ra_8_8;
  wire       [0:0]    _zz_sbuf_ra_8_9;
  wire       [0:0]    _zz_sbuf_ra_9;
  wire       [2:0]    _zz_sbuf_ra_9_1;
  wire       [3:0]    _zz_sbuf_ra_9_2;
  wire       [0:0]    _zz_sbuf_ra_9_3;
  wire       [2:0]    _zz_sbuf_ra_9_4;
  wire       [3:0]    _zz_sbuf_ra_9_5;
  wire       [0:0]    _zz_sbuf_ra_9_6;
  wire       [1:0]    _zz_sbuf_ra_9_7;
  wire       [0:0]    _zz_sbuf_ra_9_8;
  wire       [0:0]    _zz_sbuf_ra_9_9;
  wire       [0:0]    _zz_sbuf_ra_10;
  wire       [2:0]    _zz_sbuf_ra_10_1;
  wire       [3:0]    _zz_sbuf_ra_10_2;
  wire       [0:0]    _zz_sbuf_ra_10_3;
  wire       [2:0]    _zz_sbuf_ra_10_4;
  wire       [3:0]    _zz_sbuf_ra_10_5;
  wire       [0:0]    _zz_sbuf_ra_10_6;
  wire       [1:0]    _zz_sbuf_ra_10_7;
  wire       [0:0]    _zz_sbuf_ra_10_8;
  wire       [0:0]    _zz_sbuf_ra_10_9;
  wire       [0:0]    _zz_sbuf_ra_11;
  wire       [2:0]    _zz_sbuf_ra_11_1;
  wire       [3:0]    _zz_sbuf_ra_11_2;
  wire       [0:0]    _zz_sbuf_ra_11_3;
  wire       [2:0]    _zz_sbuf_ra_11_4;
  wire       [3:0]    _zz_sbuf_ra_11_5;
  wire       [0:0]    _zz_sbuf_ra_11_6;
  wire       [1:0]    _zz_sbuf_ra_11_7;
  wire       [0:0]    _zz_sbuf_ra_11_8;
  wire       [0:0]    _zz_sbuf_ra_11_9;
  wire       [0:0]    _zz_sbuf_ra_12;
  wire       [2:0]    _zz_sbuf_ra_12_1;
  wire       [3:0]    _zz_sbuf_ra_12_2;
  wire       [0:0]    _zz_sbuf_ra_12_3;
  wire       [2:0]    _zz_sbuf_ra_12_4;
  wire       [3:0]    _zz_sbuf_ra_12_5;
  wire       [0:0]    _zz_sbuf_ra_12_6;
  wire       [1:0]    _zz_sbuf_ra_12_7;
  wire       [0:0]    _zz_sbuf_ra_12_8;
  wire       [0:0]    _zz_sbuf_ra_12_9;
  wire       [0:0]    _zz_sbuf_ra_13;
  wire       [2:0]    _zz_sbuf_ra_13_1;
  wire       [3:0]    _zz_sbuf_ra_13_2;
  wire       [0:0]    _zz_sbuf_ra_13_3;
  wire       [2:0]    _zz_sbuf_ra_13_4;
  wire       [3:0]    _zz_sbuf_ra_13_5;
  wire       [0:0]    _zz_sbuf_ra_13_6;
  wire       [1:0]    _zz_sbuf_ra_13_7;
  wire       [0:0]    _zz_sbuf_ra_13_8;
  wire       [0:0]    _zz_sbuf_ra_13_9;
  wire       [0:0]    _zz_sbuf_ra_14;
  wire       [2:0]    _zz_sbuf_ra_14_1;
  wire       [3:0]    _zz_sbuf_ra_14_2;
  wire       [0:0]    _zz_sbuf_ra_14_3;
  wire       [2:0]    _zz_sbuf_ra_14_4;
  wire       [3:0]    _zz_sbuf_ra_14_5;
  wire       [0:0]    _zz_sbuf_ra_14_6;
  wire       [1:0]    _zz_sbuf_ra_14_7;
  wire       [0:0]    _zz_sbuf_ra_14_8;
  wire       [0:0]    _zz_sbuf_ra_14_9;
  wire       [0:0]    _zz_sbuf_ra_15;
  wire       [2:0]    _zz_sbuf_ra_15_1;
  wire       [3:0]    _zz_sbuf_ra_15_2;
  wire       [0:0]    _zz_sbuf_ra_15_3;
  wire       [2:0]    _zz_sbuf_ra_15_4;
  wire       [3:0]    _zz_sbuf_ra_15_5;
  wire       [0:0]    _zz_sbuf_ra_15_6;
  wire       [1:0]    _zz_sbuf_ra_15_7;
  wire       [0:0]    _zz_sbuf_ra_15_8;
  wire       [0:0]    _zz_sbuf_ra_15_9;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_1;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_2;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_3;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_4;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_5;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_6;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_7;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_8;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_9;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_10;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_11;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_12;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_13;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_14;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_15;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_16;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_17;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_18;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_19;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_20;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_21;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_22;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_23;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_24;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_25;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_26;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_27;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_28;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_29;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_30;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_31;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_32;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_33;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_34;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_35;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_36;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_37;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_38;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_39;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_40;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_41;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_42;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_43;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_44;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_45;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_46;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_47;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_48;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_49;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_50;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_51;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_52;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_53;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_54;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_55;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_56;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_57;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_58;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_59;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_60;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_61;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_62;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_63;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_64;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_65;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_66;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_67;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_68;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_69;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_70;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_71;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_72;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_73;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_74;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_75;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_76;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_77;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_78;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_79;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_80;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_81;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_82;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_83;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_84;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_85;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_86;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_87;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_88;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_89;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_90;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_91;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_92;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_93;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_94;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_95;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_96;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_97;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_98;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_99;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_100;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_101;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_102;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_103;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_104;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_105;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_106;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_107;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_108;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_109;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_110;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_111;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_112;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_113;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_114;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_115;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_116;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_117;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_118;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_119;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_120;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_121;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_122;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_123;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_124;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_125;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_126;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_127;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_128;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_129;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_130;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_131;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_132;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_133;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_134;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_135;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_136;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_137;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_138;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_139;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_140;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_141;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_142;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_143;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_144;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_145;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_146;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_147;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_148;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_149;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_150;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_151;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_152;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_153;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_154;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_155;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_156;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_157;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_158;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_159;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_160;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_161;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_162;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_163;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_164;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_165;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_166;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_167;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_168;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_169;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_170;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_171;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_172;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_173;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_174;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_175;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_176;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_177;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_178;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_179;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_180;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_181;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_182;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_183;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_184;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_185;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_186;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_187;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_188;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_189;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_190;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_191;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_192;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_193;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_194;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_195;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_196;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_197;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_198;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_199;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_200;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_201;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_202;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_203;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_204;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_205;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_206;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_207;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_208;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_209;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_210;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_211;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_212;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_213;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_214;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_215;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_216;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_217;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_218;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_219;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_220;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_221;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_222;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_223;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_224;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_225;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_226;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_227;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_228;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_229;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_230;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_231;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_232;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_233;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_234;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_235;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_236;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_237;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_238;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_239;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_240;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_241;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_242;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_243;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_244;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_245;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_246;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_247;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_248;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_249;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_250;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_251;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_252;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_253;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_254;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_255;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_256;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_257;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_258;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_259;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_260;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_261;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_262;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_263;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_264;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_265;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_266;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_267;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_268;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_269;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_270;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_271;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_272;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_273;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_274;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_275;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_276;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_277;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_278;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_279;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_280;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_281;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_282;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_283;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_284;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_285;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_286;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_287;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_288;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_289;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_290;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_291;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_292;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_293;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_294;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_295;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_296;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_297;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_298;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_299;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_300;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_301;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_302;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_303;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_304;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_305;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_306;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_307;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_308;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_309;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_310;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_311;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_312;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_313;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_314;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_315;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_316;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_317;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_318;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_319;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_320;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_321;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_322;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_323;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_324;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_325;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_326;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_327;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_328;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_329;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_330;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_331;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_332;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_333;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_334;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_335;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_336;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_337;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_338;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_339;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_340;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_341;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_342;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_343;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_344;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_345;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_346;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_347;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_348;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_349;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_350;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_351;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_352;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_353;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_354;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_355;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_356;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_357;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_358;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_359;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_360;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_361;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_362;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_363;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_364;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_365;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_366;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_367;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_368;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_369;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_370;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_371;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_372;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_373;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_374;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_375;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_376;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_377;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_378;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_379;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_380;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_381;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_382;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_383;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_384;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_385;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_386;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_387;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_388;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_389;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_390;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_391;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_392;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_393;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_394;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_395;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_396;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_397;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_398;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_399;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_400;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_401;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_402;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_403;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_404;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_405;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_406;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_407;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_408;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_409;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_410;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_411;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_412;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_413;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_414;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_415;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_416;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_417;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_418;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_419;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_420;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_421;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_422;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_423;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_424;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_425;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_426;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_427;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_428;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_429;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_430;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_431;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_432;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_433;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_434;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_435;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_436;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_437;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_438;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_439;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_440;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_441;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_442;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_443;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_444;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_445;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_446;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_447;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_448;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_449;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_450;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_451;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_452;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_453;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_454;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_455;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_456;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_457;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_458;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_459;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_460;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_461;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_462;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_463;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_464;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_465;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_466;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_467;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_468;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_469;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_470;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_471;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_472;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_473;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_474;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_475;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_476;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_477;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_478;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_479;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_480;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_481;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_482;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_483;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_484;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_485;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_486;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_487;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_488;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_489;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_490;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_491;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_492;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_493;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_494;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_495;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_496;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_497;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_498;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_499;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_500;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_501;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_502;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_503;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_504;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_505;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_506;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_507;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_508;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_509;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_510;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_511;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_512;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_513;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_514;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_515;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_516;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_517;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_518;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_519;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_520;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_521;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_522;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_523;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_524;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_525;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_526;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_527;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_528;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_529;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_530;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_531;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_532;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_533;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_534;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_535;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_536;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_537;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_538;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_539;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_540;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_541;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_542;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_543;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_544;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_545;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_546;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_547;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_548;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_549;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_550;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_551;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_552;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_553;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_554;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_555;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_556;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_557;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_558;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_559;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_560;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_561;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_562;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_563;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_564;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_565;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_566;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_567;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_568;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_569;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_570;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_571;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_572;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_573;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_574;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_575;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_576;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_577;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_578;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_579;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_580;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_581;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_582;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_583;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_584;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_585;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_586;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_587;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_588;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_589;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_590;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_591;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_592;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_593;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_594;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_595;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_596;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_597;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_598;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_599;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_600;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_601;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_602;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_603;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_604;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_605;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_606;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_607;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_608;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_609;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_610;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_611;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_612;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_613;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_614;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_615;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_616;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_617;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_618;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_619;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_620;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_621;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_622;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_623;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_624;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_625;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_626;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_627;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_628;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_629;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_630;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_631;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_632;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_633;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_634;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_635;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_636;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_637;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_638;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_639;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_640;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_641;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_642;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_643;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_644;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_645;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_646;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_647;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_648;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_649;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_650;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_651;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_652;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_653;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_654;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_655;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_656;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_657;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_658;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_659;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_660;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_661;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_662;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_663;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_664;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_665;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_666;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_667;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_668;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_669;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_670;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_671;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_672;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_673;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_674;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_675;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_676;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_677;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_678;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_679;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_680;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_681;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_682;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_683;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_684;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_685;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_686;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_687;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_688;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_689;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_690;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_691;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_692;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_693;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_694;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_695;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_696;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_697;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_698;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_699;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_700;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_701;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_702;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_703;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_704;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_705;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_706;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_707;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_708;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_709;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_710;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_711;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_712;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_713;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_714;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_715;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_716;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_717;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_718;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_719;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_720;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_721;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_722;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_723;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_724;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_725;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_726;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_727;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_728;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_729;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_730;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_731;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_732;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_733;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_734;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_735;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_736;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_737;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_738;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_739;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_740;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_741;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_742;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_743;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_744;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_745;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_746;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_747;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_748;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_749;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_750;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_751;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_752;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_753;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_754;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_755;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_756;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_757;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_758;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_759;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_760;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_761;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_762;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_763;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_764;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_765;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_766;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_767;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_768;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_769;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_770;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_771;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_772;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_773;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_774;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_775;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_776;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_777;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_778;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_779;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_780;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_781;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_782;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_783;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_784;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_785;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_786;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_787;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_788;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_789;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_790;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_791;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_792;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_793;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_794;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_795;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_796;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_797;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_798;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_799;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_800;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_801;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_802;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_803;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_804;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_805;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_806;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_807;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_808;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_809;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_810;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_811;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_812;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_813;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_814;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_815;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_816;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_817;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_818;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_819;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_820;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_821;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_822;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_823;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_824;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_825;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_826;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_827;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_828;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_829;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_830;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_831;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_832;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_833;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_834;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_835;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_836;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_837;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_838;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_839;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_840;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_841;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_842;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_843;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_844;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_845;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_846;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_847;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_848;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_849;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_850;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_851;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_852;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_853;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_854;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_855;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_856;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_857;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_858;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_859;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_860;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_861;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_862;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_863;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_864;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_865;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_866;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_867;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_868;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_869;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_870;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_871;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_872;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_873;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_874;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_875;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_876;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_877;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_878;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_879;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_880;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_881;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_882;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_883;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_884;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_885;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_886;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_887;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_888;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_889;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_890;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_891;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_892;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_893;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_894;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_895;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_896;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_897;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_898;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_899;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_900;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_901;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_902;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_903;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_904;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_905;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_906;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_907;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_908;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_909;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_910;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_911;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_912;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_913;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_914;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_915;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_916;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_917;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_918;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_919;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_920;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_921;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_922;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_923;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_924;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_925;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_926;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_927;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_928;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_929;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_930;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_931;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_932;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_933;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_934;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_935;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_936;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_937;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_938;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_939;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_940;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_941;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_942;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_943;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_944;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_945;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_946;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_947;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_948;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_949;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_950;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_951;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_952;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_953;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_954;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_955;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_956;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_957;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_958;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_959;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_960;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_961;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_962;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_963;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_964;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_965;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_966;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_967;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_968;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_969;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_970;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_971;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_972;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_973;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_974;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_975;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_976;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_977;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_978;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_979;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_980;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_981;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_982;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_983;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_984;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_985;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_986;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_987;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_988;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_989;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_990;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_991;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_992;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_993;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_994;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_995;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_996;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_997;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_998;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_999;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1000;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1001;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1002;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1003;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1004;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1005;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1006;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_1007;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_1008;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1009;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_1010;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1011;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_1012;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1013;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_1014;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1015;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_1016;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1017;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_1018;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1019;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_1020;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1021;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_1022;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1023;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1024;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1025;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1026;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1027;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1028;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1029;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1030;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1031;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1032;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1033;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1034;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1035;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1036;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1037;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1038;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1039;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1040;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1041;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1042;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1043;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1044;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1045;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1046;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1047;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1048;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1049;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1050;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1051;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1052;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1053;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1054;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1055;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1056;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1057;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1058;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1059;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1060;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1061;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1062;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1063;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1064;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1065;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1066;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1067;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1068;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1069;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1070;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1071;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1072;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1073;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1074;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1075;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1076;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1077;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1078;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1079;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1080;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1081;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1082;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1083;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1084;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1085;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1086;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1087;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1088;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1089;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1090;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1091;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1092;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1093;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1094;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1095;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1096;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1097;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1098;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1099;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1100;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1101;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1102;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1103;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1104;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1105;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1106;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1107;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1108;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1109;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1110;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1111;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1112;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1113;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1114;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1115;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1116;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1117;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_1118;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1119;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1120;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1121;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_1122;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1123;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_1124;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1125;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_1126;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1127;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_1128;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1129;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_1130;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1131;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_1132;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1133;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_1134;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1135;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1136;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1137;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1138;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1139;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1140;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1141;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1142;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1143;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1144;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1145;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1146;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1147;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1148;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1149;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1150;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1151;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1152;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1153;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1154;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1155;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1156;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1157;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1158;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1159;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1160;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1161;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1162;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1163;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1164;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1165;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1166;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1167;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1168;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1169;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1170;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1171;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1172;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1173;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1174;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1175;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1176;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1177;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1178;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1179;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1180;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1181;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1182;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1183;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1184;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1185;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1186;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1187;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1188;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1189;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1190;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1191;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1192;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1193;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1194;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1195;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1196;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1197;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1198;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1199;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1200;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1201;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1202;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1203;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1204;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1205;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1206;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1207;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1208;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1209;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1210;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1211;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1212;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1213;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1214;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1215;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1216;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1217;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1218;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1219;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1220;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1221;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1222;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1223;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1224;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1225;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1226;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1227;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1228;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1229;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1230;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1231;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_1232;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_1233;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1234;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_1235;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1236;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_1237;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1238;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_1239;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1240;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_1241;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1242;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_1243;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1244;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_1245;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1246;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1247;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1248;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1249;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1250;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1251;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1252;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1253;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1254;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1255;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1256;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1257;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1258;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1259;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1260;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1261;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1262;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1263;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1264;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1265;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1266;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1267;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1268;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1269;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1270;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1271;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1272;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1273;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1274;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1275;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1276;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1277;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1278;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1279;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1280;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1281;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1282;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1283;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1284;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1285;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1286;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1287;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1288;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1289;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1290;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1291;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1292;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1293;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1294;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1295;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1296;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1297;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1298;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1299;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1300;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1301;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1302;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1303;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1304;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1305;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1306;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1307;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1308;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1309;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1310;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1311;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1312;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1313;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1314;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1315;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1316;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1317;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1318;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1319;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1320;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1321;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1322;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1323;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1324;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1325;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1326;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1327;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1328;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1329;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1330;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1331;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1332;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1333;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1334;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1335;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1336;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1337;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1338;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1339;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1340;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1341;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1342;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_1343;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1344;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1345;
  wire       [63:0]   _zz_shareBuffer_sbuf_p0_rdat_1346;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1347;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_1348;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1349;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_1350;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1351;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_1352;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1353;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_1354;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1355;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_1356;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1357;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1358;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1359;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1360;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1361;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1362;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1363;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1364;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1365;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1366;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1367;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1368;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1369;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1370;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1371;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1372;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1373;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1374;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1375;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1376;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1377;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1378;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1379;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1380;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1381;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1382;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1383;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1384;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1385;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1386;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1387;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1388;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1389;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1390;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1391;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1392;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1393;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1394;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1395;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1396;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1397;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1398;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1399;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1400;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1401;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1402;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1403;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1404;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1405;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1406;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1407;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1408;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1409;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1410;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1411;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1412;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1413;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1414;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1415;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1416;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1417;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1418;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1419;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1420;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1421;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1422;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1423;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1424;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1425;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1426;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1427;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1428;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1429;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1430;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1431;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1432;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1433;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1434;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1435;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1436;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1437;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1438;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1439;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1440;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1441;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1442;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1443;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1444;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1445;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1446;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1447;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1448;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1449;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1450;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1451;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1452;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1453;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1454;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1455;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_1456;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1457;
  wire       [62:0]   _zz_shareBuffer_sbuf_p0_rdat_1458;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1459;
  wire       [59:0]   _zz_shareBuffer_sbuf_p0_rdat_1460;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1461;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_1462;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1463;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_1464;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1465;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_1466;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1467;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1468;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1469;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1470;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1471;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1472;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1473;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1474;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1475;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1476;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1477;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1478;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1479;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1480;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1481;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1482;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1483;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1484;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1485;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1486;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1487;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1488;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1489;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1490;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1491;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1492;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1493;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1494;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1495;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1496;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1497;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1498;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1499;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1500;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1501;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1502;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1503;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1504;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1505;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1506;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1507;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1508;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1509;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1510;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1511;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1512;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1513;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1514;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1515;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1516;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1517;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1518;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1519;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1520;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1521;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1522;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1523;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1524;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1525;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1526;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1527;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1528;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1529;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1530;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1531;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1532;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1533;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1534;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1535;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1536;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1537;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1538;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1539;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1540;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1541;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1542;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1543;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1544;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1545;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1546;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1547;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1548;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1549;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1550;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1551;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1552;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1553;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1554;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1555;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1556;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1557;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1558;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1559;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1560;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1561;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1562;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1563;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1564;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1565;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_1566;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1567;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1568;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1569;
  wire       [61:0]   _zz_shareBuffer_sbuf_p0_rdat_1570;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1571;
  wire       [58:0]   _zz_shareBuffer_sbuf_p0_rdat_1572;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1573;
  wire       [56:0]   _zz_shareBuffer_sbuf_p0_rdat_1574;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1575;
  wire       [54:0]   _zz_shareBuffer_sbuf_p0_rdat_1576;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1577;
  wire       [52:0]   _zz_shareBuffer_sbuf_p0_rdat_1578;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1579;
  wire       [50:0]   _zz_shareBuffer_sbuf_p0_rdat_1580;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1581;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1582;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1583;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1584;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1585;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1586;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1587;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1588;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1589;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1590;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1591;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1592;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1593;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1594;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1595;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1596;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1597;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1598;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1599;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1600;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1601;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1602;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1603;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1604;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1605;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1606;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1607;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1608;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1609;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1610;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1611;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1612;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1613;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1614;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1615;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1616;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1617;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1618;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1619;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1620;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1621;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1622;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1623;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1624;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1625;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1626;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1627;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1628;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1629;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1630;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1631;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1632;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1633;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1634;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1635;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1636;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1637;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1638;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1639;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1640;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1641;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1642;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1643;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1644;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1645;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1646;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1647;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1648;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1649;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1650;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1651;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1652;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1653;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1654;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1655;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1656;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1657;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1658;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1659;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1660;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1661;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1662;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1663;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1664;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1665;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1666;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1667;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1668;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1669;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1670;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1671;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1672;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1673;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1674;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1675;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_1676;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1677;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_1678;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1679;
  wire       [60:0]   _zz_shareBuffer_sbuf_p0_rdat_1680;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1681;
  wire       [57:0]   _zz_shareBuffer_sbuf_p0_rdat_1682;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1683;
  wire       [55:0]   _zz_shareBuffer_sbuf_p0_rdat_1684;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1685;
  wire       [53:0]   _zz_shareBuffer_sbuf_p0_rdat_1686;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1687;
  wire       [51:0]   _zz_shareBuffer_sbuf_p0_rdat_1688;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1689;
  wire       [49:0]   _zz_shareBuffer_sbuf_p0_rdat_1690;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1691;
  wire       [48:0]   _zz_shareBuffer_sbuf_p0_rdat_1692;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1693;
  wire       [47:0]   _zz_shareBuffer_sbuf_p0_rdat_1694;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1695;
  wire       [46:0]   _zz_shareBuffer_sbuf_p0_rdat_1696;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1697;
  wire       [45:0]   _zz_shareBuffer_sbuf_p0_rdat_1698;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1699;
  wire       [44:0]   _zz_shareBuffer_sbuf_p0_rdat_1700;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1701;
  wire       [43:0]   _zz_shareBuffer_sbuf_p0_rdat_1702;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1703;
  wire       [42:0]   _zz_shareBuffer_sbuf_p0_rdat_1704;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1705;
  wire       [41:0]   _zz_shareBuffer_sbuf_p0_rdat_1706;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1707;
  wire       [40:0]   _zz_shareBuffer_sbuf_p0_rdat_1708;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1709;
  wire       [39:0]   _zz_shareBuffer_sbuf_p0_rdat_1710;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1711;
  wire       [38:0]   _zz_shareBuffer_sbuf_p0_rdat_1712;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1713;
  wire       [37:0]   _zz_shareBuffer_sbuf_p0_rdat_1714;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1715;
  wire       [36:0]   _zz_shareBuffer_sbuf_p0_rdat_1716;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1717;
  wire       [35:0]   _zz_shareBuffer_sbuf_p0_rdat_1718;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1719;
  wire       [34:0]   _zz_shareBuffer_sbuf_p0_rdat_1720;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1721;
  wire       [33:0]   _zz_shareBuffer_sbuf_p0_rdat_1722;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1723;
  wire       [32:0]   _zz_shareBuffer_sbuf_p0_rdat_1724;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1725;
  wire       [31:0]   _zz_shareBuffer_sbuf_p0_rdat_1726;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1727;
  wire       [30:0]   _zz_shareBuffer_sbuf_p0_rdat_1728;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1729;
  wire       [29:0]   _zz_shareBuffer_sbuf_p0_rdat_1730;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1731;
  wire       [28:0]   _zz_shareBuffer_sbuf_p0_rdat_1732;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1733;
  wire       [27:0]   _zz_shareBuffer_sbuf_p0_rdat_1734;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1735;
  wire       [26:0]   _zz_shareBuffer_sbuf_p0_rdat_1736;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1737;
  wire       [25:0]   _zz_shareBuffer_sbuf_p0_rdat_1738;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1739;
  wire       [24:0]   _zz_shareBuffer_sbuf_p0_rdat_1740;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1741;
  wire       [23:0]   _zz_shareBuffer_sbuf_p0_rdat_1742;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1743;
  wire       [22:0]   _zz_shareBuffer_sbuf_p0_rdat_1744;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1745;
  wire       [21:0]   _zz_shareBuffer_sbuf_p0_rdat_1746;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1747;
  wire       [20:0]   _zz_shareBuffer_sbuf_p0_rdat_1748;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1749;
  wire       [19:0]   _zz_shareBuffer_sbuf_p0_rdat_1750;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1751;
  wire       [18:0]   _zz_shareBuffer_sbuf_p0_rdat_1752;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1753;
  wire       [17:0]   _zz_shareBuffer_sbuf_p0_rdat_1754;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1755;
  wire       [16:0]   _zz_shareBuffer_sbuf_p0_rdat_1756;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1757;
  wire       [15:0]   _zz_shareBuffer_sbuf_p0_rdat_1758;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1759;
  wire       [14:0]   _zz_shareBuffer_sbuf_p0_rdat_1760;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1761;
  wire       [13:0]   _zz_shareBuffer_sbuf_p0_rdat_1762;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1763;
  wire       [12:0]   _zz_shareBuffer_sbuf_p0_rdat_1764;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1765;
  wire       [11:0]   _zz_shareBuffer_sbuf_p0_rdat_1766;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1767;
  wire       [10:0]   _zz_shareBuffer_sbuf_p0_rdat_1768;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1769;
  wire       [9:0]    _zz_shareBuffer_sbuf_p0_rdat_1770;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1771;
  wire       [8:0]    _zz_shareBuffer_sbuf_p0_rdat_1772;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1773;
  wire       [7:0]    _zz_shareBuffer_sbuf_p0_rdat_1774;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1775;
  wire       [6:0]    _zz_shareBuffer_sbuf_p0_rdat_1776;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1777;
  wire       [5:0]    _zz_shareBuffer_sbuf_p0_rdat_1778;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1779;
  wire       [4:0]    _zz_shareBuffer_sbuf_p0_rdat_1780;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1781;
  wire       [3:0]    _zz_shareBuffer_sbuf_p0_rdat_1782;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1783;
  wire       [2:0]    _zz_shareBuffer_sbuf_p0_rdat_1784;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1785;
  wire       [1:0]    _zz_shareBuffer_sbuf_p0_rdat_1786;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1787;
  wire       [0:0]    _zz_shareBuffer_sbuf_p0_rdat_1788;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_1;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_2;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_3;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_4;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_5;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_6;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_7;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_8;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_9;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_10;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_11;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_12;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_13;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_14;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_15;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_16;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_17;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_18;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_19;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_20;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_21;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_22;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_23;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_24;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_25;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_26;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_27;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_28;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_29;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_30;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_31;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_32;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_33;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_34;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_35;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_36;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_37;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_38;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_39;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_40;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_41;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_42;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_43;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_44;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_45;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_46;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_47;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_48;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_49;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_50;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_51;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_52;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_53;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_54;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_55;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_56;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_57;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_58;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_59;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_60;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_61;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_62;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_63;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_64;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_65;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_66;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_67;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_68;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_69;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_70;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_71;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_72;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_73;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_74;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_75;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_76;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_77;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_78;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_79;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_80;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_81;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_82;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_83;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_84;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_85;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_86;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_87;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_88;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_89;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_90;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_91;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_92;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_93;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_94;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_95;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_96;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_97;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_98;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_99;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_100;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_101;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_102;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_103;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_104;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_105;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_106;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_107;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_108;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_109;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_110;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_111;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_112;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_113;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_114;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_115;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_116;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_117;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_118;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_119;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_120;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_121;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_122;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_123;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_124;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_125;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_126;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_127;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_128;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_129;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_130;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_131;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_132;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_133;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_134;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_135;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_136;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_137;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_138;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_139;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_140;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_141;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_142;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_143;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_144;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_145;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_146;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_147;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_148;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_149;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_150;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_151;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_152;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_153;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_154;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_155;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_156;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_157;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_158;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_159;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_160;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_161;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_162;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_163;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_164;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_165;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_166;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_167;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_168;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_169;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_170;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_171;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_172;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_173;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_174;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_175;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_176;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_177;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_178;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_179;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_180;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_181;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_182;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_183;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_184;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_185;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_186;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_187;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_188;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_189;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_190;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_191;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_192;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_193;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_194;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_195;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_196;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_197;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_198;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_199;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_200;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_201;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_202;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_203;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_204;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_205;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_206;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_207;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_208;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_209;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_210;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_211;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_212;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_213;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_214;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_215;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_216;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_217;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_218;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_219;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_220;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_221;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_222;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_223;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_224;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_225;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_226;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_227;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_228;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_229;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_230;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_231;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_232;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_233;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_234;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_235;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_236;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_237;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_238;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_239;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_240;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_241;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_242;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_243;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_244;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_245;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_246;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_247;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_248;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_249;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_250;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_251;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_252;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_253;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_254;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_255;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_256;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_257;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_258;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_259;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_260;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_261;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_262;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_263;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_264;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_265;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_266;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_267;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_268;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_269;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_270;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_271;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_272;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_273;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_274;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_275;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_276;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_277;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_278;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_279;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_280;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_281;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_282;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_283;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_284;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_285;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_286;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_287;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_288;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_289;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_290;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_291;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_292;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_293;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_294;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_295;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_296;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_297;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_298;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_299;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_300;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_301;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_302;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_303;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_304;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_305;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_306;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_307;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_308;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_309;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_310;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_311;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_312;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_313;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_314;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_315;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_316;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_317;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_318;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_319;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_320;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_321;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_322;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_323;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_324;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_325;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_326;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_327;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_328;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_329;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_330;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_331;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_332;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_333;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_334;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_335;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_336;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_337;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_338;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_339;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_340;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_341;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_342;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_343;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_344;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_345;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_346;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_347;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_348;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_349;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_350;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_351;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_352;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_353;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_354;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_355;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_356;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_357;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_358;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_359;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_360;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_361;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_362;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_363;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_364;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_365;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_366;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_367;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_368;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_369;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_370;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_371;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_372;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_373;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_374;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_375;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_376;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_377;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_378;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_379;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_380;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_381;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_382;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_383;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_384;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_385;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_386;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_387;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_388;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_389;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_390;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_391;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_392;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_393;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_394;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_395;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_396;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_397;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_398;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_399;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_400;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_401;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_402;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_403;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_404;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_405;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_406;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_407;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_408;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_409;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_410;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_411;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_412;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_413;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_414;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_415;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_416;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_417;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_418;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_419;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_420;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_421;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_422;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_423;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_424;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_425;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_426;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_427;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_428;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_429;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_430;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_431;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_432;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_433;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_434;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_435;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_436;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_437;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_438;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_439;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_440;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_441;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_442;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_443;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_444;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_445;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_446;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_447;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_448;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_449;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_450;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_451;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_452;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_453;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_454;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_455;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_456;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_457;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_458;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_459;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_460;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_461;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_462;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_463;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_464;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_465;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_466;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_467;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_468;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_469;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_470;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_471;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_472;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_473;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_474;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_475;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_476;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_477;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_478;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_479;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_480;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_481;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_482;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_483;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_484;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_485;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_486;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_487;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_488;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_489;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_490;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_491;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_492;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_493;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_494;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_495;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_496;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_497;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_498;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_499;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_500;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_501;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_502;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_503;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_504;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_505;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_506;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_507;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_508;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_509;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_510;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_511;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_512;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_513;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_514;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_515;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_516;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_517;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_518;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_519;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_520;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_521;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_522;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_523;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_524;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_525;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_526;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_527;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_528;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_529;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_530;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_531;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_532;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_533;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_534;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_535;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_536;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_537;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_538;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_539;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_540;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_541;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_542;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_543;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_544;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_545;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_546;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_547;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_548;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_549;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_550;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_551;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_552;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_553;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_554;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_555;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_556;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_557;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_558;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_559;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_560;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_561;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_562;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_563;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_564;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_565;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_566;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_567;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_568;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_569;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_570;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_571;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_572;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_573;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_574;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_575;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_576;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_577;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_578;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_579;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_580;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_581;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_582;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_583;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_584;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_585;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_586;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_587;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_588;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_589;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_590;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_591;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_592;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_593;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_594;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_595;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_596;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_597;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_598;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_599;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_600;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_601;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_602;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_603;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_604;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_605;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_606;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_607;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_608;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_609;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_610;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_611;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_612;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_613;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_614;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_615;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_616;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_617;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_618;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_619;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_620;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_621;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_622;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_623;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_624;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_625;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_626;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_627;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_628;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_629;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_630;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_631;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_632;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_633;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_634;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_635;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_636;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_637;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_638;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_639;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_640;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_641;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_642;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_643;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_644;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_645;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_646;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_647;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_648;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_649;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_650;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_651;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_652;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_653;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_654;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_655;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_656;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_657;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_658;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_659;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_660;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_661;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_662;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_663;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_664;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_665;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_666;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_667;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_668;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_669;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_670;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_671;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_672;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_673;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_674;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_675;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_676;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_677;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_678;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_679;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_680;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_681;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_682;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_683;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_684;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_685;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_686;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_687;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_688;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_689;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_690;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_691;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_692;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_693;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_694;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_695;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_696;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_697;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_698;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_699;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_700;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_701;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_702;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_703;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_704;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_705;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_706;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_707;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_708;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_709;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_710;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_711;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_712;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_713;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_714;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_715;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_716;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_717;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_718;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_719;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_720;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_721;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_722;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_723;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_724;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_725;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_726;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_727;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_728;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_729;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_730;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_731;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_732;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_733;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_734;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_735;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_736;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_737;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_738;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_739;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_740;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_741;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_742;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_743;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_744;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_745;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_746;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_747;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_748;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_749;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_750;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_751;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_752;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_753;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_754;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_755;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_756;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_757;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_758;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_759;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_760;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_761;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_762;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_763;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_764;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_765;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_766;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_767;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_768;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_769;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_770;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_771;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_772;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_773;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_774;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_775;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_776;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_777;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_778;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_779;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_780;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_781;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_782;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_783;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_784;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_785;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_786;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_787;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_788;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_789;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_790;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_791;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_792;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_793;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_794;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_795;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_796;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_797;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_798;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_799;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_800;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_801;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_802;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_803;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_804;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_805;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_806;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_807;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_808;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_809;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_810;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_811;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_812;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_813;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_814;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_815;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_816;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_817;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_818;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_819;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_820;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_821;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_822;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_823;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_824;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_825;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_826;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_827;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_828;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_829;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_830;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_831;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_832;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_833;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_834;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_835;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_836;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_837;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_838;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_839;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_840;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_841;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_842;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_843;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_844;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_845;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_846;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_847;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_848;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_849;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_850;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_851;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_852;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_853;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_854;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_855;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_856;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_857;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_858;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_859;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_860;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_861;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_862;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_863;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_864;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_865;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_866;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_867;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_868;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_869;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_870;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_871;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_872;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_873;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_874;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_875;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_876;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_877;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_878;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_879;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_880;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_881;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_882;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_883;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_884;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_885;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_886;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_887;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_888;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_889;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_890;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_891;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_892;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_893;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_894;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_895;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_896;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_897;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_898;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_899;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_900;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_901;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_902;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_903;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_904;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_905;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_906;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_907;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_908;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_909;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_910;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_911;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_912;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_913;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_914;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_915;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_916;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_917;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_918;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_919;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_920;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_921;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_922;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_923;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_924;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_925;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_926;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_927;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_928;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_929;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_930;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_931;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_932;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_933;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_934;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_935;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_936;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_937;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_938;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_939;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_940;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_941;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_942;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_943;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_944;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_945;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_946;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_947;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_948;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_949;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_950;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_951;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_952;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_953;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_954;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_955;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_956;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_957;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_958;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_959;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_960;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_961;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_962;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_963;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_964;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_965;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_966;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_967;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_968;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_969;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_970;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_971;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_972;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_973;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_974;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_975;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_976;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_977;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_978;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_979;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_980;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_981;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_982;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_983;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_984;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_985;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_986;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_987;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_988;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_989;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_990;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_991;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_992;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_993;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_994;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_995;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_996;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_997;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_998;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_999;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1000;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1001;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1002;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1003;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1004;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1005;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1006;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_1007;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_1008;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1009;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_1010;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1011;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_1012;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1013;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_1014;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1015;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_1016;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1017;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_1018;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1019;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_1020;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1021;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_1022;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1023;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1024;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1025;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1026;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1027;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1028;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1029;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1030;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1031;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1032;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1033;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1034;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1035;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1036;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1037;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1038;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1039;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1040;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1041;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1042;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1043;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1044;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1045;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1046;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1047;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1048;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1049;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1050;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1051;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1052;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1053;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1054;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1055;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1056;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1057;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1058;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1059;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1060;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1061;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1062;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1063;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1064;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1065;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1066;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1067;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1068;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1069;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1070;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1071;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1072;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1073;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1074;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1075;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1076;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1077;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1078;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1079;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1080;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1081;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1082;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1083;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1084;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1085;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1086;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1087;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1088;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1089;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1090;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1091;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1092;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1093;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1094;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1095;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1096;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1097;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1098;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1099;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1100;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1101;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1102;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1103;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1104;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1105;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1106;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1107;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1108;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1109;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1110;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1111;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1112;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1113;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1114;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1115;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1116;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1117;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_1118;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1119;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1120;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1121;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_1122;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1123;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_1124;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1125;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_1126;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1127;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_1128;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1129;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_1130;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1131;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_1132;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1133;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_1134;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1135;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1136;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1137;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1138;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1139;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1140;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1141;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1142;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1143;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1144;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1145;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1146;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1147;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1148;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1149;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1150;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1151;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1152;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1153;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1154;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1155;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1156;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1157;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1158;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1159;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1160;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1161;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1162;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1163;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1164;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1165;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1166;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1167;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1168;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1169;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1170;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1171;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1172;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1173;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1174;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1175;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1176;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1177;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1178;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1179;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1180;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1181;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1182;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1183;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1184;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1185;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1186;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1187;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1188;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1189;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1190;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1191;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1192;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1193;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1194;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1195;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1196;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1197;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1198;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1199;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1200;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1201;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1202;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1203;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1204;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1205;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1206;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1207;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1208;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1209;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1210;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1211;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1212;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1213;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1214;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1215;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1216;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1217;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1218;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1219;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1220;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1221;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1222;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1223;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1224;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1225;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1226;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1227;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1228;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1229;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1230;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1231;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_1232;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_1233;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1234;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_1235;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1236;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_1237;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1238;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_1239;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1240;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_1241;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1242;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_1243;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1244;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_1245;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1246;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1247;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1248;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1249;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1250;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1251;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1252;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1253;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1254;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1255;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1256;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1257;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1258;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1259;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1260;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1261;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1262;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1263;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1264;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1265;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1266;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1267;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1268;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1269;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1270;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1271;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1272;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1273;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1274;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1275;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1276;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1277;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1278;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1279;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1280;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1281;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1282;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1283;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1284;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1285;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1286;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1287;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1288;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1289;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1290;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1291;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1292;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1293;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1294;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1295;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1296;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1297;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1298;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1299;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1300;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1301;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1302;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1303;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1304;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1305;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1306;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1307;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1308;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1309;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1310;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1311;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1312;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1313;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1314;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1315;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1316;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1317;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1318;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1319;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1320;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1321;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1322;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1323;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1324;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1325;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1326;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1327;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1328;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1329;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1330;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1331;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1332;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1333;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1334;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1335;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1336;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1337;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1338;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1339;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1340;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1341;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1342;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_1343;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1344;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1345;
  wire       [63:0]   _zz_shareBuffer_sbuf_p1_rdat_1346;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1347;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_1348;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1349;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_1350;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1351;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_1352;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1353;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_1354;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1355;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_1356;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1357;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1358;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1359;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1360;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1361;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1362;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1363;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1364;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1365;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1366;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1367;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1368;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1369;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1370;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1371;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1372;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1373;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1374;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1375;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1376;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1377;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1378;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1379;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1380;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1381;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1382;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1383;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1384;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1385;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1386;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1387;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1388;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1389;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1390;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1391;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1392;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1393;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1394;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1395;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1396;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1397;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1398;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1399;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1400;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1401;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1402;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1403;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1404;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1405;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1406;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1407;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1408;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1409;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1410;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1411;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1412;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1413;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1414;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1415;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1416;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1417;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1418;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1419;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1420;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1421;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1422;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1423;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1424;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1425;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1426;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1427;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1428;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1429;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1430;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1431;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1432;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1433;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1434;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1435;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1436;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1437;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1438;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1439;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1440;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1441;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1442;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1443;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1444;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1445;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1446;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1447;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1448;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1449;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1450;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1451;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1452;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1453;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1454;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1455;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_1456;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1457;
  wire       [62:0]   _zz_shareBuffer_sbuf_p1_rdat_1458;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1459;
  wire       [59:0]   _zz_shareBuffer_sbuf_p1_rdat_1460;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1461;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_1462;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1463;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_1464;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1465;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_1466;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1467;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1468;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1469;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1470;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1471;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1472;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1473;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1474;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1475;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1476;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1477;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1478;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1479;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1480;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1481;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1482;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1483;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1484;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1485;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1486;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1487;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1488;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1489;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1490;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1491;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1492;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1493;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1494;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1495;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1496;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1497;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1498;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1499;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1500;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1501;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1502;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1503;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1504;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1505;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1506;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1507;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1508;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1509;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1510;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1511;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1512;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1513;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1514;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1515;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1516;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1517;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1518;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1519;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1520;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1521;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1522;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1523;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1524;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1525;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1526;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1527;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1528;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1529;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1530;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1531;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1532;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1533;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1534;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1535;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1536;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1537;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1538;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1539;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1540;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1541;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1542;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1543;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1544;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1545;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1546;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1547;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1548;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1549;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1550;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1551;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1552;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1553;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1554;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1555;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1556;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1557;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1558;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1559;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1560;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1561;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1562;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1563;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1564;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1565;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_1566;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1567;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1568;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1569;
  wire       [61:0]   _zz_shareBuffer_sbuf_p1_rdat_1570;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1571;
  wire       [58:0]   _zz_shareBuffer_sbuf_p1_rdat_1572;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1573;
  wire       [56:0]   _zz_shareBuffer_sbuf_p1_rdat_1574;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1575;
  wire       [54:0]   _zz_shareBuffer_sbuf_p1_rdat_1576;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1577;
  wire       [52:0]   _zz_shareBuffer_sbuf_p1_rdat_1578;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1579;
  wire       [50:0]   _zz_shareBuffer_sbuf_p1_rdat_1580;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1581;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1582;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1583;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1584;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1585;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1586;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1587;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1588;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1589;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1590;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1591;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1592;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1593;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1594;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1595;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1596;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1597;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1598;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1599;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1600;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1601;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1602;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1603;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1604;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1605;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1606;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1607;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1608;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1609;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1610;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1611;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1612;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1613;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1614;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1615;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1616;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1617;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1618;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1619;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1620;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1621;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1622;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1623;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1624;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1625;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1626;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1627;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1628;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1629;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1630;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1631;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1632;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1633;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1634;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1635;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1636;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1637;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1638;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1639;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1640;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1641;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1642;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1643;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1644;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1645;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1646;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1647;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1648;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1649;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1650;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1651;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1652;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1653;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1654;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1655;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1656;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1657;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1658;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1659;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1660;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1661;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1662;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1663;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1664;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1665;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1666;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1667;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1668;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1669;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1670;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1671;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1672;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1673;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1674;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1675;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_1676;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1677;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_1678;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1679;
  wire       [60:0]   _zz_shareBuffer_sbuf_p1_rdat_1680;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1681;
  wire       [57:0]   _zz_shareBuffer_sbuf_p1_rdat_1682;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1683;
  wire       [55:0]   _zz_shareBuffer_sbuf_p1_rdat_1684;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1685;
  wire       [53:0]   _zz_shareBuffer_sbuf_p1_rdat_1686;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1687;
  wire       [51:0]   _zz_shareBuffer_sbuf_p1_rdat_1688;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1689;
  wire       [49:0]   _zz_shareBuffer_sbuf_p1_rdat_1690;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1691;
  wire       [48:0]   _zz_shareBuffer_sbuf_p1_rdat_1692;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1693;
  wire       [47:0]   _zz_shareBuffer_sbuf_p1_rdat_1694;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1695;
  wire       [46:0]   _zz_shareBuffer_sbuf_p1_rdat_1696;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1697;
  wire       [45:0]   _zz_shareBuffer_sbuf_p1_rdat_1698;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1699;
  wire       [44:0]   _zz_shareBuffer_sbuf_p1_rdat_1700;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1701;
  wire       [43:0]   _zz_shareBuffer_sbuf_p1_rdat_1702;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1703;
  wire       [42:0]   _zz_shareBuffer_sbuf_p1_rdat_1704;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1705;
  wire       [41:0]   _zz_shareBuffer_sbuf_p1_rdat_1706;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1707;
  wire       [40:0]   _zz_shareBuffer_sbuf_p1_rdat_1708;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1709;
  wire       [39:0]   _zz_shareBuffer_sbuf_p1_rdat_1710;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1711;
  wire       [38:0]   _zz_shareBuffer_sbuf_p1_rdat_1712;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1713;
  wire       [37:0]   _zz_shareBuffer_sbuf_p1_rdat_1714;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1715;
  wire       [36:0]   _zz_shareBuffer_sbuf_p1_rdat_1716;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1717;
  wire       [35:0]   _zz_shareBuffer_sbuf_p1_rdat_1718;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1719;
  wire       [34:0]   _zz_shareBuffer_sbuf_p1_rdat_1720;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1721;
  wire       [33:0]   _zz_shareBuffer_sbuf_p1_rdat_1722;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1723;
  wire       [32:0]   _zz_shareBuffer_sbuf_p1_rdat_1724;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1725;
  wire       [31:0]   _zz_shareBuffer_sbuf_p1_rdat_1726;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1727;
  wire       [30:0]   _zz_shareBuffer_sbuf_p1_rdat_1728;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1729;
  wire       [29:0]   _zz_shareBuffer_sbuf_p1_rdat_1730;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1731;
  wire       [28:0]   _zz_shareBuffer_sbuf_p1_rdat_1732;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1733;
  wire       [27:0]   _zz_shareBuffer_sbuf_p1_rdat_1734;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1735;
  wire       [26:0]   _zz_shareBuffer_sbuf_p1_rdat_1736;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1737;
  wire       [25:0]   _zz_shareBuffer_sbuf_p1_rdat_1738;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1739;
  wire       [24:0]   _zz_shareBuffer_sbuf_p1_rdat_1740;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1741;
  wire       [23:0]   _zz_shareBuffer_sbuf_p1_rdat_1742;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1743;
  wire       [22:0]   _zz_shareBuffer_sbuf_p1_rdat_1744;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1745;
  wire       [21:0]   _zz_shareBuffer_sbuf_p1_rdat_1746;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1747;
  wire       [20:0]   _zz_shareBuffer_sbuf_p1_rdat_1748;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1749;
  wire       [19:0]   _zz_shareBuffer_sbuf_p1_rdat_1750;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1751;
  wire       [18:0]   _zz_shareBuffer_sbuf_p1_rdat_1752;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1753;
  wire       [17:0]   _zz_shareBuffer_sbuf_p1_rdat_1754;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1755;
  wire       [16:0]   _zz_shareBuffer_sbuf_p1_rdat_1756;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1757;
  wire       [15:0]   _zz_shareBuffer_sbuf_p1_rdat_1758;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1759;
  wire       [14:0]   _zz_shareBuffer_sbuf_p1_rdat_1760;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1761;
  wire       [13:0]   _zz_shareBuffer_sbuf_p1_rdat_1762;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1763;
  wire       [12:0]   _zz_shareBuffer_sbuf_p1_rdat_1764;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1765;
  wire       [11:0]   _zz_shareBuffer_sbuf_p1_rdat_1766;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1767;
  wire       [10:0]   _zz_shareBuffer_sbuf_p1_rdat_1768;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1769;
  wire       [9:0]    _zz_shareBuffer_sbuf_p1_rdat_1770;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1771;
  wire       [8:0]    _zz_shareBuffer_sbuf_p1_rdat_1772;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1773;
  wire       [7:0]    _zz_shareBuffer_sbuf_p1_rdat_1774;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1775;
  wire       [6:0]    _zz_shareBuffer_sbuf_p1_rdat_1776;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1777;
  wire       [5:0]    _zz_shareBuffer_sbuf_p1_rdat_1778;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1779;
  wire       [4:0]    _zz_shareBuffer_sbuf_p1_rdat_1780;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1781;
  wire       [3:0]    _zz_shareBuffer_sbuf_p1_rdat_1782;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1783;
  wire       [2:0]    _zz_shareBuffer_sbuf_p1_rdat_1784;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1785;
  wire       [1:0]    _zz_shareBuffer_sbuf_p1_rdat_1786;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1787;
  wire       [0:0]    _zz_shareBuffer_sbuf_p1_rdat_1788;
  wire       [3:0]    dc2sbuf_p0_wr_bsel;
  wire       [3:0]    img2sbuf_p0_wr_bsel;
  wire       [3:0]    dc2sbuf_p1_wr_bsel;
  wire       [3:0]    img2sbuf_p1_wr_bsel;
  wire                dc2sbuf_p0_wr_sel_0;
  wire                dc2sbuf_p0_wr_sel_1;
  wire                dc2sbuf_p0_wr_sel_2;
  wire                dc2sbuf_p0_wr_sel_3;
  wire                dc2sbuf_p0_wr_sel_4;
  wire                dc2sbuf_p0_wr_sel_5;
  wire                dc2sbuf_p0_wr_sel_6;
  wire                dc2sbuf_p0_wr_sel_7;
  wire                dc2sbuf_p0_wr_sel_8;
  wire                dc2sbuf_p0_wr_sel_9;
  wire                dc2sbuf_p0_wr_sel_10;
  wire                dc2sbuf_p0_wr_sel_11;
  wire                dc2sbuf_p0_wr_sel_12;
  wire                dc2sbuf_p0_wr_sel_13;
  wire                dc2sbuf_p0_wr_sel_14;
  wire                dc2sbuf_p0_wr_sel_15;
  wire                dc2sbuf_p1_wr_sel_0;
  wire                dc2sbuf_p1_wr_sel_1;
  wire                dc2sbuf_p1_wr_sel_2;
  wire                dc2sbuf_p1_wr_sel_3;
  wire                dc2sbuf_p1_wr_sel_4;
  wire                dc2sbuf_p1_wr_sel_5;
  wire                dc2sbuf_p1_wr_sel_6;
  wire                dc2sbuf_p1_wr_sel_7;
  wire                dc2sbuf_p1_wr_sel_8;
  wire                dc2sbuf_p1_wr_sel_9;
  wire                dc2sbuf_p1_wr_sel_10;
  wire                dc2sbuf_p1_wr_sel_11;
  wire                dc2sbuf_p1_wr_sel_12;
  wire                dc2sbuf_p1_wr_sel_13;
  wire                dc2sbuf_p1_wr_sel_14;
  wire                dc2sbuf_p1_wr_sel_15;
  wire                img2sbuf_p0_wr_sel_0;
  wire                img2sbuf_p0_wr_sel_1;
  wire                img2sbuf_p0_wr_sel_2;
  wire                img2sbuf_p0_wr_sel_3;
  wire                img2sbuf_p0_wr_sel_4;
  wire                img2sbuf_p0_wr_sel_5;
  wire                img2sbuf_p0_wr_sel_6;
  wire                img2sbuf_p0_wr_sel_7;
  wire                img2sbuf_p0_wr_sel_8;
  wire                img2sbuf_p0_wr_sel_9;
  wire                img2sbuf_p0_wr_sel_10;
  wire                img2sbuf_p0_wr_sel_11;
  wire                img2sbuf_p0_wr_sel_12;
  wire                img2sbuf_p0_wr_sel_13;
  wire                img2sbuf_p0_wr_sel_14;
  wire                img2sbuf_p0_wr_sel_15;
  wire                img2sbuf_p1_wr_sel_0;
  wire                img2sbuf_p1_wr_sel_1;
  wire                img2sbuf_p1_wr_sel_2;
  wire                img2sbuf_p1_wr_sel_3;
  wire                img2sbuf_p1_wr_sel_4;
  wire                img2sbuf_p1_wr_sel_5;
  wire                img2sbuf_p1_wr_sel_6;
  wire                img2sbuf_p1_wr_sel_7;
  wire                img2sbuf_p1_wr_sel_8;
  wire                img2sbuf_p1_wr_sel_9;
  wire                img2sbuf_p1_wr_sel_10;
  wire                img2sbuf_p1_wr_sel_11;
  wire                img2sbuf_p1_wr_sel_12;
  wire                img2sbuf_p1_wr_sel_13;
  wire                img2sbuf_p1_wr_sel_14;
  wire                img2sbuf_p1_wr_sel_15;
  wire                sbuf_we_0;
  wire                sbuf_we_1;
  wire                sbuf_we_2;
  wire                sbuf_we_3;
  wire                sbuf_we_4;
  wire                sbuf_we_5;
  wire                sbuf_we_6;
  wire                sbuf_we_7;
  wire                sbuf_we_8;
  wire                sbuf_we_9;
  wire                sbuf_we_10;
  wire                sbuf_we_11;
  wire                sbuf_we_12;
  wire                sbuf_we_13;
  wire                sbuf_we_14;
  wire                sbuf_we_15;
  wire       [3:0]    sbuf_wa_0;
  wire       [3:0]    sbuf_wa_1;
  wire       [3:0]    sbuf_wa_2;
  wire       [3:0]    sbuf_wa_3;
  wire       [3:0]    sbuf_wa_4;
  wire       [3:0]    sbuf_wa_5;
  wire       [3:0]    sbuf_wa_6;
  wire       [3:0]    sbuf_wa_7;
  wire       [3:0]    sbuf_wa_8;
  wire       [3:0]    sbuf_wa_9;
  wire       [3:0]    sbuf_wa_10;
  wire       [3:0]    sbuf_wa_11;
  wire       [3:0]    sbuf_wa_12;
  wire       [3:0]    sbuf_wa_13;
  wire       [3:0]    sbuf_wa_14;
  wire       [3:0]    sbuf_wa_15;
  wire       [63:0]   sbuf_wdat_0;
  wire       [63:0]   sbuf_wdat_1;
  wire       [63:0]   sbuf_wdat_2;
  wire       [63:0]   sbuf_wdat_3;
  wire       [63:0]   sbuf_wdat_4;
  wire       [63:0]   sbuf_wdat_5;
  wire       [63:0]   sbuf_wdat_6;
  wire       [63:0]   sbuf_wdat_7;
  wire       [63:0]   sbuf_wdat_8;
  wire       [63:0]   sbuf_wdat_9;
  wire       [63:0]   sbuf_wdat_10;
  wire       [63:0]   sbuf_wdat_11;
  wire       [63:0]   sbuf_wdat_12;
  wire       [63:0]   sbuf_wdat_13;
  wire       [63:0]   sbuf_wdat_14;
  wire       [63:0]   sbuf_wdat_15;
  wire       [3:0]    dc2sbuf_p0_rd_bsel;
  wire       [3:0]    img2sbuf_p0_rd_bsel;
  wire       [3:0]    dc2sbuf_p1_rd_bsel;
  wire       [3:0]    img2sbuf_p1_rd_bsel;
  wire                dc2sbuf_p0_rd_sel_0;
  wire                dc2sbuf_p0_rd_sel_1;
  wire                dc2sbuf_p0_rd_sel_2;
  wire                dc2sbuf_p0_rd_sel_3;
  wire                dc2sbuf_p0_rd_sel_4;
  wire                dc2sbuf_p0_rd_sel_5;
  wire                dc2sbuf_p0_rd_sel_6;
  wire                dc2sbuf_p0_rd_sel_7;
  wire                dc2sbuf_p0_rd_sel_8;
  wire                dc2sbuf_p0_rd_sel_9;
  wire                dc2sbuf_p0_rd_sel_10;
  wire                dc2sbuf_p0_rd_sel_11;
  wire                dc2sbuf_p0_rd_sel_12;
  wire                dc2sbuf_p0_rd_sel_13;
  wire                dc2sbuf_p0_rd_sel_14;
  wire                dc2sbuf_p0_rd_sel_15;
  wire                dc2sbuf_p1_rd_sel_0;
  wire                dc2sbuf_p1_rd_sel_1;
  wire                dc2sbuf_p1_rd_sel_2;
  wire                dc2sbuf_p1_rd_sel_3;
  wire                dc2sbuf_p1_rd_sel_4;
  wire                dc2sbuf_p1_rd_sel_5;
  wire                dc2sbuf_p1_rd_sel_6;
  wire                dc2sbuf_p1_rd_sel_7;
  wire                dc2sbuf_p1_rd_sel_8;
  wire                dc2sbuf_p1_rd_sel_9;
  wire                dc2sbuf_p1_rd_sel_10;
  wire                dc2sbuf_p1_rd_sel_11;
  wire                dc2sbuf_p1_rd_sel_12;
  wire                dc2sbuf_p1_rd_sel_13;
  wire                dc2sbuf_p1_rd_sel_14;
  wire                dc2sbuf_p1_rd_sel_15;
  wire                img2sbuf_p0_rd_sel_0;
  wire                img2sbuf_p0_rd_sel_1;
  wire                img2sbuf_p0_rd_sel_2;
  wire                img2sbuf_p0_rd_sel_3;
  wire                img2sbuf_p0_rd_sel_4;
  wire                img2sbuf_p0_rd_sel_5;
  wire                img2sbuf_p0_rd_sel_6;
  wire                img2sbuf_p0_rd_sel_7;
  wire                img2sbuf_p0_rd_sel_8;
  wire                img2sbuf_p0_rd_sel_9;
  wire                img2sbuf_p0_rd_sel_10;
  wire                img2sbuf_p0_rd_sel_11;
  wire                img2sbuf_p0_rd_sel_12;
  wire                img2sbuf_p0_rd_sel_13;
  wire                img2sbuf_p0_rd_sel_14;
  wire                img2sbuf_p0_rd_sel_15;
  wire                img2sbuf_p1_rd_sel_0;
  wire                img2sbuf_p1_rd_sel_1;
  wire                img2sbuf_p1_rd_sel_2;
  wire                img2sbuf_p1_rd_sel_3;
  wire                img2sbuf_p1_rd_sel_4;
  wire                img2sbuf_p1_rd_sel_5;
  wire                img2sbuf_p1_rd_sel_6;
  wire                img2sbuf_p1_rd_sel_7;
  wire                img2sbuf_p1_rd_sel_8;
  wire                img2sbuf_p1_rd_sel_9;
  wire                img2sbuf_p1_rd_sel_10;
  wire                img2sbuf_p1_rd_sel_11;
  wire                img2sbuf_p1_rd_sel_12;
  wire                img2sbuf_p1_rd_sel_13;
  wire                img2sbuf_p1_rd_sel_14;
  wire                img2sbuf_p1_rd_sel_15;
  wire                sbuf_p0_re_0;
  wire                sbuf_p0_re_1;
  wire                sbuf_p0_re_2;
  wire                sbuf_p0_re_3;
  wire                sbuf_p0_re_4;
  wire                sbuf_p0_re_5;
  wire                sbuf_p0_re_6;
  wire                sbuf_p0_re_7;
  wire                sbuf_p0_re_8;
  wire                sbuf_p0_re_9;
  wire                sbuf_p0_re_10;
  wire                sbuf_p0_re_11;
  wire                sbuf_p0_re_12;
  wire                sbuf_p0_re_13;
  wire                sbuf_p0_re_14;
  wire                sbuf_p0_re_15;
  wire                sbuf_p1_re_0;
  wire                sbuf_p1_re_1;
  wire                sbuf_p1_re_2;
  wire                sbuf_p1_re_3;
  wire                sbuf_p1_re_4;
  wire                sbuf_p1_re_5;
  wire                sbuf_p1_re_6;
  wire                sbuf_p1_re_7;
  wire                sbuf_p1_re_8;
  wire                sbuf_p1_re_9;
  wire                sbuf_p1_re_10;
  wire                sbuf_p1_re_11;
  wire                sbuf_p1_re_12;
  wire                sbuf_p1_re_13;
  wire                sbuf_p1_re_14;
  wire                sbuf_p1_re_15;
  wire                sbuf_re_0;
  wire                sbuf_re_1;
  wire                sbuf_re_2;
  wire                sbuf_re_3;
  wire                sbuf_re_4;
  wire                sbuf_re_5;
  wire                sbuf_re_6;
  wire                sbuf_re_7;
  wire                sbuf_re_8;
  wire                sbuf_re_9;
  wire                sbuf_re_10;
  wire                sbuf_re_11;
  wire                sbuf_re_12;
  wire                sbuf_re_13;
  wire                sbuf_re_14;
  wire                sbuf_re_15;
  wire       [3:0]    sbuf_ra_0;
  wire       [3:0]    sbuf_ra_1;
  wire       [3:0]    sbuf_ra_2;
  wire       [3:0]    sbuf_ra_3;
  wire       [3:0]    sbuf_ra_4;
  wire       [3:0]    sbuf_ra_5;
  wire       [3:0]    sbuf_ra_6;
  wire       [3:0]    sbuf_ra_7;
  wire       [3:0]    sbuf_ra_8;
  wire       [3:0]    sbuf_ra_9;
  wire       [3:0]    sbuf_ra_10;
  wire       [3:0]    sbuf_ra_11;
  wire       [3:0]    sbuf_ra_12;
  wire       [3:0]    sbuf_ra_13;
  wire       [3:0]    sbuf_ra_14;
  wire       [3:0]    sbuf_ra_15;
  wire       [63:0]   shareBuffer_sbuf_rdat_0;
  wire       [63:0]   shareBuffer_sbuf_rdat_1;
  wire       [63:0]   shareBuffer_sbuf_rdat_2;
  wire       [63:0]   shareBuffer_sbuf_rdat_3;
  wire       [63:0]   shareBuffer_sbuf_rdat_4;
  wire       [63:0]   shareBuffer_sbuf_rdat_5;
  wire       [63:0]   shareBuffer_sbuf_rdat_6;
  wire       [63:0]   shareBuffer_sbuf_rdat_7;
  wire       [63:0]   shareBuffer_sbuf_rdat_8;
  wire       [63:0]   shareBuffer_sbuf_rdat_9;
  wire       [63:0]   shareBuffer_sbuf_rdat_10;
  wire       [63:0]   shareBuffer_sbuf_rdat_11;
  wire       [63:0]   shareBuffer_sbuf_rdat_12;
  wire       [63:0]   shareBuffer_sbuf_rdat_13;
  wire       [63:0]   shareBuffer_sbuf_rdat_14;
  wire       [63:0]   shareBuffer_sbuf_rdat_15;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_0;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_1;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_2;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_3;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_4;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_5;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_6;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_7;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_8;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_9;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_10;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_11;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_12;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_13;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_14;
  reg                 shareBuffer_sbuf_p0_re_norm_d1_15;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_0;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_1;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_2;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_3;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_4;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_5;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_6;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_7;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_8;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_9;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_10;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_11;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_12;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_13;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_14;
  reg                 shareBuffer_sbuf_p1_re_norm_d1_15;
  reg                 shareBuffer_sbuf_p0_rd_en_d1;
  reg                 shareBuffer_sbuf_p1_rd_en_d1;
  wire       [63:0]   shareBuffer_sbuf_p0_rdat;
  wire       [63:0]   shareBuffer_sbuf_p1_rdat;
  reg        [63:0]   shareBuffer_sbuf_p0_rdat_d2;
  reg        [63:0]   shareBuffer_sbuf_p1_rdat_d2;

  assign _zz_sbuf_wa_0 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wa_0_1 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,dc2sbuf_p0_wr_sel_0}};
  assign _zz_sbuf_wa_0_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_0_3 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wa_0_4 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,dc2sbuf_p1_wr_sel_0}};
  assign _zz_sbuf_wa_0_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_0_6 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wa_0_7 = {img2sbuf_p0_wr_sel_0,img2sbuf_p0_wr_sel_0};
  assign _zz_sbuf_wa_0_8 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wa_0_9 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wa_1 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wa_1_1 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,dc2sbuf_p0_wr_sel_1}};
  assign _zz_sbuf_wa_1_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_1_3 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wa_1_4 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,dc2sbuf_p1_wr_sel_1}};
  assign _zz_sbuf_wa_1_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_1_6 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wa_1_7 = {img2sbuf_p0_wr_sel_1,img2sbuf_p0_wr_sel_1};
  assign _zz_sbuf_wa_1_8 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wa_1_9 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wa_2 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wa_2_1 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,dc2sbuf_p0_wr_sel_2}};
  assign _zz_sbuf_wa_2_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_2_3 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wa_2_4 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,dc2sbuf_p1_wr_sel_2}};
  assign _zz_sbuf_wa_2_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_2_6 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wa_2_7 = {img2sbuf_p0_wr_sel_2,img2sbuf_p0_wr_sel_2};
  assign _zz_sbuf_wa_2_8 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wa_2_9 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wa_3 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wa_3_1 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,dc2sbuf_p0_wr_sel_3}};
  assign _zz_sbuf_wa_3_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_3_3 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wa_3_4 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,dc2sbuf_p1_wr_sel_3}};
  assign _zz_sbuf_wa_3_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_3_6 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wa_3_7 = {img2sbuf_p0_wr_sel_3,img2sbuf_p0_wr_sel_3};
  assign _zz_sbuf_wa_3_8 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wa_3_9 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wa_4 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wa_4_1 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,dc2sbuf_p0_wr_sel_4}};
  assign _zz_sbuf_wa_4_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_4_3 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wa_4_4 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,dc2sbuf_p1_wr_sel_4}};
  assign _zz_sbuf_wa_4_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_4_6 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wa_4_7 = {img2sbuf_p0_wr_sel_4,img2sbuf_p0_wr_sel_4};
  assign _zz_sbuf_wa_4_8 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wa_4_9 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wa_5 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wa_5_1 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,dc2sbuf_p0_wr_sel_5}};
  assign _zz_sbuf_wa_5_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_5_3 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wa_5_4 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,dc2sbuf_p1_wr_sel_5}};
  assign _zz_sbuf_wa_5_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_5_6 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wa_5_7 = {img2sbuf_p0_wr_sel_5,img2sbuf_p0_wr_sel_5};
  assign _zz_sbuf_wa_5_8 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wa_5_9 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wa_6 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wa_6_1 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,dc2sbuf_p0_wr_sel_6}};
  assign _zz_sbuf_wa_6_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_6_3 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wa_6_4 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,dc2sbuf_p1_wr_sel_6}};
  assign _zz_sbuf_wa_6_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_6_6 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wa_6_7 = {img2sbuf_p0_wr_sel_6,img2sbuf_p0_wr_sel_6};
  assign _zz_sbuf_wa_6_8 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wa_6_9 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wa_7 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wa_7_1 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,dc2sbuf_p0_wr_sel_7}};
  assign _zz_sbuf_wa_7_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_7_3 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wa_7_4 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,dc2sbuf_p1_wr_sel_7}};
  assign _zz_sbuf_wa_7_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_7_6 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wa_7_7 = {img2sbuf_p0_wr_sel_7,img2sbuf_p0_wr_sel_7};
  assign _zz_sbuf_wa_7_8 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wa_7_9 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wa_8 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wa_8_1 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,dc2sbuf_p0_wr_sel_8}};
  assign _zz_sbuf_wa_8_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_8_3 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wa_8_4 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,dc2sbuf_p1_wr_sel_8}};
  assign _zz_sbuf_wa_8_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_8_6 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wa_8_7 = {img2sbuf_p0_wr_sel_8,img2sbuf_p0_wr_sel_8};
  assign _zz_sbuf_wa_8_8 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wa_8_9 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wa_9 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wa_9_1 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,dc2sbuf_p0_wr_sel_9}};
  assign _zz_sbuf_wa_9_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_9_3 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wa_9_4 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,dc2sbuf_p1_wr_sel_9}};
  assign _zz_sbuf_wa_9_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_9_6 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wa_9_7 = {img2sbuf_p0_wr_sel_9,img2sbuf_p0_wr_sel_9};
  assign _zz_sbuf_wa_9_8 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wa_9_9 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wa_10 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wa_10_1 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,dc2sbuf_p0_wr_sel_10}};
  assign _zz_sbuf_wa_10_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_10_3 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wa_10_4 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,dc2sbuf_p1_wr_sel_10}};
  assign _zz_sbuf_wa_10_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_10_6 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wa_10_7 = {img2sbuf_p0_wr_sel_10,img2sbuf_p0_wr_sel_10};
  assign _zz_sbuf_wa_10_8 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wa_10_9 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wa_11 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wa_11_1 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,dc2sbuf_p0_wr_sel_11}};
  assign _zz_sbuf_wa_11_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_11_3 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wa_11_4 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,dc2sbuf_p1_wr_sel_11}};
  assign _zz_sbuf_wa_11_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_11_6 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wa_11_7 = {img2sbuf_p0_wr_sel_11,img2sbuf_p0_wr_sel_11};
  assign _zz_sbuf_wa_11_8 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wa_11_9 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wa_12 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wa_12_1 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,dc2sbuf_p0_wr_sel_12}};
  assign _zz_sbuf_wa_12_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_12_3 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wa_12_4 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,dc2sbuf_p1_wr_sel_12}};
  assign _zz_sbuf_wa_12_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_12_6 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wa_12_7 = {img2sbuf_p0_wr_sel_12,img2sbuf_p0_wr_sel_12};
  assign _zz_sbuf_wa_12_8 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wa_12_9 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wa_13 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wa_13_1 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,dc2sbuf_p0_wr_sel_13}};
  assign _zz_sbuf_wa_13_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_13_3 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wa_13_4 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,dc2sbuf_p1_wr_sel_13}};
  assign _zz_sbuf_wa_13_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_13_6 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wa_13_7 = {img2sbuf_p0_wr_sel_13,img2sbuf_p0_wr_sel_13};
  assign _zz_sbuf_wa_13_8 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wa_13_9 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wa_14 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wa_14_1 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,dc2sbuf_p0_wr_sel_14}};
  assign _zz_sbuf_wa_14_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_14_3 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wa_14_4 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,dc2sbuf_p1_wr_sel_14}};
  assign _zz_sbuf_wa_14_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_14_6 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wa_14_7 = {img2sbuf_p0_wr_sel_14,img2sbuf_p0_wr_sel_14};
  assign _zz_sbuf_wa_14_8 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wa_14_9 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wa_15 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wa_15_1 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,dc2sbuf_p0_wr_sel_15}};
  assign _zz_sbuf_wa_15_2 = dc2sbuf_p_wr_0_addr_payload[3 : 0];
  assign _zz_sbuf_wa_15_3 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wa_15_4 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,dc2sbuf_p1_wr_sel_15}};
  assign _zz_sbuf_wa_15_5 = dc2sbuf_p_wr_1_addr_payload[3 : 0];
  assign _zz_sbuf_wa_15_6 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wa_15_7 = {img2sbuf_p0_wr_sel_15,img2sbuf_p0_wr_sel_15};
  assign _zz_sbuf_wa_15_8 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wa_15_9 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_0 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_1 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_2,_zz_sbuf_wdat_0_3}}}};
  assign _zz_sbuf_wdat_0_32 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_33 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_34,_zz_sbuf_wdat_0_35}}}};
  assign _zz_sbuf_wdat_0_64 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_65 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_66,_zz_sbuf_wdat_0_67}}}};
  assign _zz_sbuf_wdat_0_94 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_95 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_96,_zz_sbuf_wdat_0_97}}}};
  assign _zz_sbuf_wdat_0_2 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_3 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_4,_zz_sbuf_wdat_0_5}}}};
  assign _zz_sbuf_wdat_0_34 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_35 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_36,_zz_sbuf_wdat_0_37}}}};
  assign _zz_sbuf_wdat_0_66 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_67 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_68,_zz_sbuf_wdat_0_69}}}};
  assign _zz_sbuf_wdat_0_96 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_97 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_98,_zz_sbuf_wdat_0_99}}}};
  assign _zz_sbuf_wdat_0_4 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_5 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_6,_zz_sbuf_wdat_0_7}}}};
  assign _zz_sbuf_wdat_0_36 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_37 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_38,_zz_sbuf_wdat_0_39}}}};
  assign _zz_sbuf_wdat_0_68 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_69 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_70,_zz_sbuf_wdat_0_71}}}};
  assign _zz_sbuf_wdat_0_98 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_99 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_100,_zz_sbuf_wdat_0_101}}}};
  assign _zz_sbuf_wdat_0_6 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_7 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_8,_zz_sbuf_wdat_0_9}}}};
  assign _zz_sbuf_wdat_0_38 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_39 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_40,_zz_sbuf_wdat_0_41}}}};
  assign _zz_sbuf_wdat_0_70 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_71 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_72,_zz_sbuf_wdat_0_73}}}};
  assign _zz_sbuf_wdat_0_100 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_101 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_102,_zz_sbuf_wdat_0_103}}}};
  assign _zz_sbuf_wdat_0_8 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_9 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_10,_zz_sbuf_wdat_0_11}}}};
  assign _zz_sbuf_wdat_0_40 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_41 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_42,_zz_sbuf_wdat_0_43}}}};
  assign _zz_sbuf_wdat_0_72 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_73 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_74,_zz_sbuf_wdat_0_75}}}};
  assign _zz_sbuf_wdat_0_102 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_103 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_104,_zz_sbuf_wdat_0_105}}}};
  assign _zz_sbuf_wdat_0_10 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_11 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_12,_zz_sbuf_wdat_0_13}}}};
  assign _zz_sbuf_wdat_0_42 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_43 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_44,_zz_sbuf_wdat_0_45}}}};
  assign _zz_sbuf_wdat_0_74 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_75 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_76,_zz_sbuf_wdat_0_77}}}};
  assign _zz_sbuf_wdat_0_104 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_105 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_106,_zz_sbuf_wdat_0_107}}}};
  assign _zz_sbuf_wdat_0_12 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_13 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_14,_zz_sbuf_wdat_0_15}}}};
  assign _zz_sbuf_wdat_0_44 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_45 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_46,_zz_sbuf_wdat_0_47}}}};
  assign _zz_sbuf_wdat_0_76 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_77 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_78,_zz_sbuf_wdat_0_79}}}};
  assign _zz_sbuf_wdat_0_106 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_107 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_108,_zz_sbuf_wdat_0_109}}}};
  assign _zz_sbuf_wdat_0_14 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_15 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_16,_zz_sbuf_wdat_0_17}}}};
  assign _zz_sbuf_wdat_0_46 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_47 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_48,_zz_sbuf_wdat_0_49}}}};
  assign _zz_sbuf_wdat_0_78 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_79 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_80,_zz_sbuf_wdat_0_81}}}};
  assign _zz_sbuf_wdat_0_108 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_109 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_110,_zz_sbuf_wdat_0_111}}}};
  assign _zz_sbuf_wdat_0_16 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_17 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_18,_zz_sbuf_wdat_0_19}}}};
  assign _zz_sbuf_wdat_0_48 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_49 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_50,_zz_sbuf_wdat_0_51}}}};
  assign _zz_sbuf_wdat_0_80 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_81 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_82,_zz_sbuf_wdat_0_83}}}};
  assign _zz_sbuf_wdat_0_110 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_111 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_112,_zz_sbuf_wdat_0_113}}}};
  assign _zz_sbuf_wdat_0_18 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_19 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_20,_zz_sbuf_wdat_0_21}}}};
  assign _zz_sbuf_wdat_0_50 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_51 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_52,_zz_sbuf_wdat_0_53}}}};
  assign _zz_sbuf_wdat_0_82 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_83 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_84,_zz_sbuf_wdat_0_85}}}};
  assign _zz_sbuf_wdat_0_112 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_113 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_114,_zz_sbuf_wdat_0_115}}}};
  assign _zz_sbuf_wdat_0_20 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_21 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_22,_zz_sbuf_wdat_0_23}}}};
  assign _zz_sbuf_wdat_0_52 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_53 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_54,_zz_sbuf_wdat_0_55}}}};
  assign _zz_sbuf_wdat_0_84 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_85 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_86,_zz_sbuf_wdat_0_87}}}};
  assign _zz_sbuf_wdat_0_114 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_115 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_116,_zz_sbuf_wdat_0_117}}}};
  assign _zz_sbuf_wdat_0_22 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_23 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_24,_zz_sbuf_wdat_0_25}}}};
  assign _zz_sbuf_wdat_0_54 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_55 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_56,_zz_sbuf_wdat_0_57}}}};
  assign _zz_sbuf_wdat_0_86 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_87 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_88,_zz_sbuf_wdat_0_89}}}};
  assign _zz_sbuf_wdat_0_116 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_117 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_118,_zz_sbuf_wdat_0_119}}}};
  assign _zz_sbuf_wdat_0_24 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_25 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_26,_zz_sbuf_wdat_0_27}}}};
  assign _zz_sbuf_wdat_0_56 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_57 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_58,_zz_sbuf_wdat_0_59}}}};
  assign _zz_sbuf_wdat_0_88 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_89 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_90,_zz_sbuf_wdat_0_91}}}};
  assign _zz_sbuf_wdat_0_118 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_119 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_120,_zz_sbuf_wdat_0_121}}}};
  assign _zz_sbuf_wdat_0_26 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_27 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_28,_zz_sbuf_wdat_0_29}}}};
  assign _zz_sbuf_wdat_0_58 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_59 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_60,_zz_sbuf_wdat_0_61}}}};
  assign _zz_sbuf_wdat_0_90 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_91 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_92,_zz_sbuf_wdat_0_93}}}};
  assign _zz_sbuf_wdat_0_120 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_121 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_122,_zz_sbuf_wdat_0_123}}}};
  assign _zz_sbuf_wdat_0_28 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_29 = {dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_30,_zz_sbuf_wdat_0_31}}}}};
  assign _zz_sbuf_wdat_0_60 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_61 = {dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_62,_zz_sbuf_wdat_0_63}}}}};
  assign _zz_sbuf_wdat_0_92 = img2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_93 = {img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,img2sbuf_p0_wr_sel_0}}}};
  assign _zz_sbuf_wdat_0_122 = img2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_123 = {img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,img2sbuf_p1_wr_sel_0}}};
  assign _zz_sbuf_wdat_0_30 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_31 = dc2sbuf_p0_wr_sel_0;
  assign _zz_sbuf_wdat_0_62 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_0_63 = dc2sbuf_p1_wr_sel_0;
  assign _zz_sbuf_wdat_1 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_1 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_2,_zz_sbuf_wdat_1_3}}}};
  assign _zz_sbuf_wdat_1_32 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_33 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_34,_zz_sbuf_wdat_1_35}}}};
  assign _zz_sbuf_wdat_1_64 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_65 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_66,_zz_sbuf_wdat_1_67}}}};
  assign _zz_sbuf_wdat_1_94 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_95 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_96,_zz_sbuf_wdat_1_97}}}};
  assign _zz_sbuf_wdat_1_2 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_3 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_4,_zz_sbuf_wdat_1_5}}}};
  assign _zz_sbuf_wdat_1_34 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_35 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_36,_zz_sbuf_wdat_1_37}}}};
  assign _zz_sbuf_wdat_1_66 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_67 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_68,_zz_sbuf_wdat_1_69}}}};
  assign _zz_sbuf_wdat_1_96 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_97 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_98,_zz_sbuf_wdat_1_99}}}};
  assign _zz_sbuf_wdat_1_4 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_5 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_6,_zz_sbuf_wdat_1_7}}}};
  assign _zz_sbuf_wdat_1_36 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_37 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_38,_zz_sbuf_wdat_1_39}}}};
  assign _zz_sbuf_wdat_1_68 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_69 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_70,_zz_sbuf_wdat_1_71}}}};
  assign _zz_sbuf_wdat_1_98 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_99 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_100,_zz_sbuf_wdat_1_101}}}};
  assign _zz_sbuf_wdat_1_6 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_7 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_8,_zz_sbuf_wdat_1_9}}}};
  assign _zz_sbuf_wdat_1_38 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_39 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_40,_zz_sbuf_wdat_1_41}}}};
  assign _zz_sbuf_wdat_1_70 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_71 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_72,_zz_sbuf_wdat_1_73}}}};
  assign _zz_sbuf_wdat_1_100 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_101 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_102,_zz_sbuf_wdat_1_103}}}};
  assign _zz_sbuf_wdat_1_8 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_9 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_10,_zz_sbuf_wdat_1_11}}}};
  assign _zz_sbuf_wdat_1_40 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_41 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_42,_zz_sbuf_wdat_1_43}}}};
  assign _zz_sbuf_wdat_1_72 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_73 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_74,_zz_sbuf_wdat_1_75}}}};
  assign _zz_sbuf_wdat_1_102 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_103 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_104,_zz_sbuf_wdat_1_105}}}};
  assign _zz_sbuf_wdat_1_10 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_11 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_12,_zz_sbuf_wdat_1_13}}}};
  assign _zz_sbuf_wdat_1_42 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_43 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_44,_zz_sbuf_wdat_1_45}}}};
  assign _zz_sbuf_wdat_1_74 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_75 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_76,_zz_sbuf_wdat_1_77}}}};
  assign _zz_sbuf_wdat_1_104 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_105 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_106,_zz_sbuf_wdat_1_107}}}};
  assign _zz_sbuf_wdat_1_12 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_13 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_14,_zz_sbuf_wdat_1_15}}}};
  assign _zz_sbuf_wdat_1_44 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_45 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_46,_zz_sbuf_wdat_1_47}}}};
  assign _zz_sbuf_wdat_1_76 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_77 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_78,_zz_sbuf_wdat_1_79}}}};
  assign _zz_sbuf_wdat_1_106 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_107 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_108,_zz_sbuf_wdat_1_109}}}};
  assign _zz_sbuf_wdat_1_14 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_15 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_16,_zz_sbuf_wdat_1_17}}}};
  assign _zz_sbuf_wdat_1_46 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_47 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_48,_zz_sbuf_wdat_1_49}}}};
  assign _zz_sbuf_wdat_1_78 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_79 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_80,_zz_sbuf_wdat_1_81}}}};
  assign _zz_sbuf_wdat_1_108 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_109 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_110,_zz_sbuf_wdat_1_111}}}};
  assign _zz_sbuf_wdat_1_16 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_17 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_18,_zz_sbuf_wdat_1_19}}}};
  assign _zz_sbuf_wdat_1_48 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_49 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_50,_zz_sbuf_wdat_1_51}}}};
  assign _zz_sbuf_wdat_1_80 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_81 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_82,_zz_sbuf_wdat_1_83}}}};
  assign _zz_sbuf_wdat_1_110 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_111 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_112,_zz_sbuf_wdat_1_113}}}};
  assign _zz_sbuf_wdat_1_18 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_19 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_20,_zz_sbuf_wdat_1_21}}}};
  assign _zz_sbuf_wdat_1_50 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_51 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_52,_zz_sbuf_wdat_1_53}}}};
  assign _zz_sbuf_wdat_1_82 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_83 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_84,_zz_sbuf_wdat_1_85}}}};
  assign _zz_sbuf_wdat_1_112 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_113 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_114,_zz_sbuf_wdat_1_115}}}};
  assign _zz_sbuf_wdat_1_20 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_21 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_22,_zz_sbuf_wdat_1_23}}}};
  assign _zz_sbuf_wdat_1_52 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_53 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_54,_zz_sbuf_wdat_1_55}}}};
  assign _zz_sbuf_wdat_1_84 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_85 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_86,_zz_sbuf_wdat_1_87}}}};
  assign _zz_sbuf_wdat_1_114 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_115 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_116,_zz_sbuf_wdat_1_117}}}};
  assign _zz_sbuf_wdat_1_22 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_23 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_24,_zz_sbuf_wdat_1_25}}}};
  assign _zz_sbuf_wdat_1_54 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_55 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_56,_zz_sbuf_wdat_1_57}}}};
  assign _zz_sbuf_wdat_1_86 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_87 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_88,_zz_sbuf_wdat_1_89}}}};
  assign _zz_sbuf_wdat_1_116 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_117 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_118,_zz_sbuf_wdat_1_119}}}};
  assign _zz_sbuf_wdat_1_24 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_25 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_26,_zz_sbuf_wdat_1_27}}}};
  assign _zz_sbuf_wdat_1_56 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_57 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_58,_zz_sbuf_wdat_1_59}}}};
  assign _zz_sbuf_wdat_1_88 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_89 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_90,_zz_sbuf_wdat_1_91}}}};
  assign _zz_sbuf_wdat_1_118 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_119 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_120,_zz_sbuf_wdat_1_121}}}};
  assign _zz_sbuf_wdat_1_26 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_27 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_28,_zz_sbuf_wdat_1_29}}}};
  assign _zz_sbuf_wdat_1_58 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_59 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_60,_zz_sbuf_wdat_1_61}}}};
  assign _zz_sbuf_wdat_1_90 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_91 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_92,_zz_sbuf_wdat_1_93}}}};
  assign _zz_sbuf_wdat_1_120 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_121 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_122,_zz_sbuf_wdat_1_123}}}};
  assign _zz_sbuf_wdat_1_28 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_29 = {dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_30,_zz_sbuf_wdat_1_31}}}}};
  assign _zz_sbuf_wdat_1_60 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_61 = {dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_62,_zz_sbuf_wdat_1_63}}}}};
  assign _zz_sbuf_wdat_1_92 = img2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_93 = {img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,img2sbuf_p0_wr_sel_1}}}};
  assign _zz_sbuf_wdat_1_122 = img2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_123 = {img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,img2sbuf_p1_wr_sel_1}}};
  assign _zz_sbuf_wdat_1_30 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_31 = dc2sbuf_p0_wr_sel_1;
  assign _zz_sbuf_wdat_1_62 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_1_63 = dc2sbuf_p1_wr_sel_1;
  assign _zz_sbuf_wdat_2 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_1 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_2,_zz_sbuf_wdat_2_3}}}};
  assign _zz_sbuf_wdat_2_32 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_33 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_34,_zz_sbuf_wdat_2_35}}}};
  assign _zz_sbuf_wdat_2_64 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_65 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_66,_zz_sbuf_wdat_2_67}}}};
  assign _zz_sbuf_wdat_2_94 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_95 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_96,_zz_sbuf_wdat_2_97}}}};
  assign _zz_sbuf_wdat_2_2 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_3 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_4,_zz_sbuf_wdat_2_5}}}};
  assign _zz_sbuf_wdat_2_34 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_35 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_36,_zz_sbuf_wdat_2_37}}}};
  assign _zz_sbuf_wdat_2_66 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_67 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_68,_zz_sbuf_wdat_2_69}}}};
  assign _zz_sbuf_wdat_2_96 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_97 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_98,_zz_sbuf_wdat_2_99}}}};
  assign _zz_sbuf_wdat_2_4 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_5 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_6,_zz_sbuf_wdat_2_7}}}};
  assign _zz_sbuf_wdat_2_36 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_37 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_38,_zz_sbuf_wdat_2_39}}}};
  assign _zz_sbuf_wdat_2_68 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_69 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_70,_zz_sbuf_wdat_2_71}}}};
  assign _zz_sbuf_wdat_2_98 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_99 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_100,_zz_sbuf_wdat_2_101}}}};
  assign _zz_sbuf_wdat_2_6 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_7 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_8,_zz_sbuf_wdat_2_9}}}};
  assign _zz_sbuf_wdat_2_38 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_39 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_40,_zz_sbuf_wdat_2_41}}}};
  assign _zz_sbuf_wdat_2_70 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_71 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_72,_zz_sbuf_wdat_2_73}}}};
  assign _zz_sbuf_wdat_2_100 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_101 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_102,_zz_sbuf_wdat_2_103}}}};
  assign _zz_sbuf_wdat_2_8 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_9 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_10,_zz_sbuf_wdat_2_11}}}};
  assign _zz_sbuf_wdat_2_40 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_41 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_42,_zz_sbuf_wdat_2_43}}}};
  assign _zz_sbuf_wdat_2_72 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_73 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_74,_zz_sbuf_wdat_2_75}}}};
  assign _zz_sbuf_wdat_2_102 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_103 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_104,_zz_sbuf_wdat_2_105}}}};
  assign _zz_sbuf_wdat_2_10 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_11 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_12,_zz_sbuf_wdat_2_13}}}};
  assign _zz_sbuf_wdat_2_42 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_43 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_44,_zz_sbuf_wdat_2_45}}}};
  assign _zz_sbuf_wdat_2_74 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_75 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_76,_zz_sbuf_wdat_2_77}}}};
  assign _zz_sbuf_wdat_2_104 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_105 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_106,_zz_sbuf_wdat_2_107}}}};
  assign _zz_sbuf_wdat_2_12 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_13 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_14,_zz_sbuf_wdat_2_15}}}};
  assign _zz_sbuf_wdat_2_44 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_45 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_46,_zz_sbuf_wdat_2_47}}}};
  assign _zz_sbuf_wdat_2_76 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_77 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_78,_zz_sbuf_wdat_2_79}}}};
  assign _zz_sbuf_wdat_2_106 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_107 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_108,_zz_sbuf_wdat_2_109}}}};
  assign _zz_sbuf_wdat_2_14 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_15 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_16,_zz_sbuf_wdat_2_17}}}};
  assign _zz_sbuf_wdat_2_46 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_47 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_48,_zz_sbuf_wdat_2_49}}}};
  assign _zz_sbuf_wdat_2_78 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_79 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_80,_zz_sbuf_wdat_2_81}}}};
  assign _zz_sbuf_wdat_2_108 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_109 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_110,_zz_sbuf_wdat_2_111}}}};
  assign _zz_sbuf_wdat_2_16 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_17 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_18,_zz_sbuf_wdat_2_19}}}};
  assign _zz_sbuf_wdat_2_48 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_49 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_50,_zz_sbuf_wdat_2_51}}}};
  assign _zz_sbuf_wdat_2_80 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_81 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_82,_zz_sbuf_wdat_2_83}}}};
  assign _zz_sbuf_wdat_2_110 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_111 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_112,_zz_sbuf_wdat_2_113}}}};
  assign _zz_sbuf_wdat_2_18 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_19 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_20,_zz_sbuf_wdat_2_21}}}};
  assign _zz_sbuf_wdat_2_50 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_51 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_52,_zz_sbuf_wdat_2_53}}}};
  assign _zz_sbuf_wdat_2_82 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_83 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_84,_zz_sbuf_wdat_2_85}}}};
  assign _zz_sbuf_wdat_2_112 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_113 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_114,_zz_sbuf_wdat_2_115}}}};
  assign _zz_sbuf_wdat_2_20 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_21 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_22,_zz_sbuf_wdat_2_23}}}};
  assign _zz_sbuf_wdat_2_52 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_53 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_54,_zz_sbuf_wdat_2_55}}}};
  assign _zz_sbuf_wdat_2_84 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_85 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_86,_zz_sbuf_wdat_2_87}}}};
  assign _zz_sbuf_wdat_2_114 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_115 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_116,_zz_sbuf_wdat_2_117}}}};
  assign _zz_sbuf_wdat_2_22 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_23 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_24,_zz_sbuf_wdat_2_25}}}};
  assign _zz_sbuf_wdat_2_54 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_55 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_56,_zz_sbuf_wdat_2_57}}}};
  assign _zz_sbuf_wdat_2_86 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_87 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_88,_zz_sbuf_wdat_2_89}}}};
  assign _zz_sbuf_wdat_2_116 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_117 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_118,_zz_sbuf_wdat_2_119}}}};
  assign _zz_sbuf_wdat_2_24 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_25 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_26,_zz_sbuf_wdat_2_27}}}};
  assign _zz_sbuf_wdat_2_56 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_57 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_58,_zz_sbuf_wdat_2_59}}}};
  assign _zz_sbuf_wdat_2_88 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_89 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_90,_zz_sbuf_wdat_2_91}}}};
  assign _zz_sbuf_wdat_2_118 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_119 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_120,_zz_sbuf_wdat_2_121}}}};
  assign _zz_sbuf_wdat_2_26 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_27 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_28,_zz_sbuf_wdat_2_29}}}};
  assign _zz_sbuf_wdat_2_58 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_59 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_60,_zz_sbuf_wdat_2_61}}}};
  assign _zz_sbuf_wdat_2_90 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_91 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_92,_zz_sbuf_wdat_2_93}}}};
  assign _zz_sbuf_wdat_2_120 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_121 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_122,_zz_sbuf_wdat_2_123}}}};
  assign _zz_sbuf_wdat_2_28 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_29 = {dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_30,_zz_sbuf_wdat_2_31}}}}};
  assign _zz_sbuf_wdat_2_60 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_61 = {dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_62,_zz_sbuf_wdat_2_63}}}}};
  assign _zz_sbuf_wdat_2_92 = img2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_93 = {img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,img2sbuf_p0_wr_sel_2}}}};
  assign _zz_sbuf_wdat_2_122 = img2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_123 = {img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,img2sbuf_p1_wr_sel_2}}};
  assign _zz_sbuf_wdat_2_30 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_31 = dc2sbuf_p0_wr_sel_2;
  assign _zz_sbuf_wdat_2_62 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_2_63 = dc2sbuf_p1_wr_sel_2;
  assign _zz_sbuf_wdat_3 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_1 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_2,_zz_sbuf_wdat_3_3}}}};
  assign _zz_sbuf_wdat_3_32 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_33 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_34,_zz_sbuf_wdat_3_35}}}};
  assign _zz_sbuf_wdat_3_64 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_65 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_66,_zz_sbuf_wdat_3_67}}}};
  assign _zz_sbuf_wdat_3_94 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_95 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_96,_zz_sbuf_wdat_3_97}}}};
  assign _zz_sbuf_wdat_3_2 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_3 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_4,_zz_sbuf_wdat_3_5}}}};
  assign _zz_sbuf_wdat_3_34 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_35 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_36,_zz_sbuf_wdat_3_37}}}};
  assign _zz_sbuf_wdat_3_66 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_67 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_68,_zz_sbuf_wdat_3_69}}}};
  assign _zz_sbuf_wdat_3_96 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_97 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_98,_zz_sbuf_wdat_3_99}}}};
  assign _zz_sbuf_wdat_3_4 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_5 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_6,_zz_sbuf_wdat_3_7}}}};
  assign _zz_sbuf_wdat_3_36 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_37 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_38,_zz_sbuf_wdat_3_39}}}};
  assign _zz_sbuf_wdat_3_68 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_69 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_70,_zz_sbuf_wdat_3_71}}}};
  assign _zz_sbuf_wdat_3_98 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_99 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_100,_zz_sbuf_wdat_3_101}}}};
  assign _zz_sbuf_wdat_3_6 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_7 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_8,_zz_sbuf_wdat_3_9}}}};
  assign _zz_sbuf_wdat_3_38 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_39 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_40,_zz_sbuf_wdat_3_41}}}};
  assign _zz_sbuf_wdat_3_70 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_71 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_72,_zz_sbuf_wdat_3_73}}}};
  assign _zz_sbuf_wdat_3_100 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_101 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_102,_zz_sbuf_wdat_3_103}}}};
  assign _zz_sbuf_wdat_3_8 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_9 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_10,_zz_sbuf_wdat_3_11}}}};
  assign _zz_sbuf_wdat_3_40 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_41 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_42,_zz_sbuf_wdat_3_43}}}};
  assign _zz_sbuf_wdat_3_72 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_73 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_74,_zz_sbuf_wdat_3_75}}}};
  assign _zz_sbuf_wdat_3_102 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_103 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_104,_zz_sbuf_wdat_3_105}}}};
  assign _zz_sbuf_wdat_3_10 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_11 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_12,_zz_sbuf_wdat_3_13}}}};
  assign _zz_sbuf_wdat_3_42 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_43 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_44,_zz_sbuf_wdat_3_45}}}};
  assign _zz_sbuf_wdat_3_74 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_75 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_76,_zz_sbuf_wdat_3_77}}}};
  assign _zz_sbuf_wdat_3_104 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_105 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_106,_zz_sbuf_wdat_3_107}}}};
  assign _zz_sbuf_wdat_3_12 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_13 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_14,_zz_sbuf_wdat_3_15}}}};
  assign _zz_sbuf_wdat_3_44 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_45 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_46,_zz_sbuf_wdat_3_47}}}};
  assign _zz_sbuf_wdat_3_76 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_77 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_78,_zz_sbuf_wdat_3_79}}}};
  assign _zz_sbuf_wdat_3_106 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_107 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_108,_zz_sbuf_wdat_3_109}}}};
  assign _zz_sbuf_wdat_3_14 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_15 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_16,_zz_sbuf_wdat_3_17}}}};
  assign _zz_sbuf_wdat_3_46 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_47 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_48,_zz_sbuf_wdat_3_49}}}};
  assign _zz_sbuf_wdat_3_78 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_79 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_80,_zz_sbuf_wdat_3_81}}}};
  assign _zz_sbuf_wdat_3_108 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_109 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_110,_zz_sbuf_wdat_3_111}}}};
  assign _zz_sbuf_wdat_3_16 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_17 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_18,_zz_sbuf_wdat_3_19}}}};
  assign _zz_sbuf_wdat_3_48 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_49 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_50,_zz_sbuf_wdat_3_51}}}};
  assign _zz_sbuf_wdat_3_80 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_81 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_82,_zz_sbuf_wdat_3_83}}}};
  assign _zz_sbuf_wdat_3_110 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_111 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_112,_zz_sbuf_wdat_3_113}}}};
  assign _zz_sbuf_wdat_3_18 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_19 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_20,_zz_sbuf_wdat_3_21}}}};
  assign _zz_sbuf_wdat_3_50 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_51 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_52,_zz_sbuf_wdat_3_53}}}};
  assign _zz_sbuf_wdat_3_82 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_83 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_84,_zz_sbuf_wdat_3_85}}}};
  assign _zz_sbuf_wdat_3_112 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_113 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_114,_zz_sbuf_wdat_3_115}}}};
  assign _zz_sbuf_wdat_3_20 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_21 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_22,_zz_sbuf_wdat_3_23}}}};
  assign _zz_sbuf_wdat_3_52 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_53 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_54,_zz_sbuf_wdat_3_55}}}};
  assign _zz_sbuf_wdat_3_84 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_85 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_86,_zz_sbuf_wdat_3_87}}}};
  assign _zz_sbuf_wdat_3_114 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_115 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_116,_zz_sbuf_wdat_3_117}}}};
  assign _zz_sbuf_wdat_3_22 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_23 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_24,_zz_sbuf_wdat_3_25}}}};
  assign _zz_sbuf_wdat_3_54 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_55 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_56,_zz_sbuf_wdat_3_57}}}};
  assign _zz_sbuf_wdat_3_86 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_87 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_88,_zz_sbuf_wdat_3_89}}}};
  assign _zz_sbuf_wdat_3_116 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_117 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_118,_zz_sbuf_wdat_3_119}}}};
  assign _zz_sbuf_wdat_3_24 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_25 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_26,_zz_sbuf_wdat_3_27}}}};
  assign _zz_sbuf_wdat_3_56 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_57 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_58,_zz_sbuf_wdat_3_59}}}};
  assign _zz_sbuf_wdat_3_88 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_89 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_90,_zz_sbuf_wdat_3_91}}}};
  assign _zz_sbuf_wdat_3_118 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_119 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_120,_zz_sbuf_wdat_3_121}}}};
  assign _zz_sbuf_wdat_3_26 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_27 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_28,_zz_sbuf_wdat_3_29}}}};
  assign _zz_sbuf_wdat_3_58 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_59 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_60,_zz_sbuf_wdat_3_61}}}};
  assign _zz_sbuf_wdat_3_90 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_91 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_92,_zz_sbuf_wdat_3_93}}}};
  assign _zz_sbuf_wdat_3_120 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_121 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_122,_zz_sbuf_wdat_3_123}}}};
  assign _zz_sbuf_wdat_3_28 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_29 = {dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_30,_zz_sbuf_wdat_3_31}}}}};
  assign _zz_sbuf_wdat_3_60 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_61 = {dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_62,_zz_sbuf_wdat_3_63}}}}};
  assign _zz_sbuf_wdat_3_92 = img2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_93 = {img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,img2sbuf_p0_wr_sel_3}}}};
  assign _zz_sbuf_wdat_3_122 = img2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_123 = {img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,img2sbuf_p1_wr_sel_3}}};
  assign _zz_sbuf_wdat_3_30 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_31 = dc2sbuf_p0_wr_sel_3;
  assign _zz_sbuf_wdat_3_62 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_3_63 = dc2sbuf_p1_wr_sel_3;
  assign _zz_sbuf_wdat_4 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_1 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_2,_zz_sbuf_wdat_4_3}}}};
  assign _zz_sbuf_wdat_4_32 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_33 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_34,_zz_sbuf_wdat_4_35}}}};
  assign _zz_sbuf_wdat_4_64 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_65 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_66,_zz_sbuf_wdat_4_67}}}};
  assign _zz_sbuf_wdat_4_94 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_95 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_96,_zz_sbuf_wdat_4_97}}}};
  assign _zz_sbuf_wdat_4_2 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_3 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_4,_zz_sbuf_wdat_4_5}}}};
  assign _zz_sbuf_wdat_4_34 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_35 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_36,_zz_sbuf_wdat_4_37}}}};
  assign _zz_sbuf_wdat_4_66 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_67 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_68,_zz_sbuf_wdat_4_69}}}};
  assign _zz_sbuf_wdat_4_96 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_97 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_98,_zz_sbuf_wdat_4_99}}}};
  assign _zz_sbuf_wdat_4_4 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_5 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_6,_zz_sbuf_wdat_4_7}}}};
  assign _zz_sbuf_wdat_4_36 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_37 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_38,_zz_sbuf_wdat_4_39}}}};
  assign _zz_sbuf_wdat_4_68 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_69 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_70,_zz_sbuf_wdat_4_71}}}};
  assign _zz_sbuf_wdat_4_98 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_99 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_100,_zz_sbuf_wdat_4_101}}}};
  assign _zz_sbuf_wdat_4_6 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_7 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_8,_zz_sbuf_wdat_4_9}}}};
  assign _zz_sbuf_wdat_4_38 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_39 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_40,_zz_sbuf_wdat_4_41}}}};
  assign _zz_sbuf_wdat_4_70 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_71 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_72,_zz_sbuf_wdat_4_73}}}};
  assign _zz_sbuf_wdat_4_100 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_101 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_102,_zz_sbuf_wdat_4_103}}}};
  assign _zz_sbuf_wdat_4_8 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_9 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_10,_zz_sbuf_wdat_4_11}}}};
  assign _zz_sbuf_wdat_4_40 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_41 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_42,_zz_sbuf_wdat_4_43}}}};
  assign _zz_sbuf_wdat_4_72 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_73 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_74,_zz_sbuf_wdat_4_75}}}};
  assign _zz_sbuf_wdat_4_102 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_103 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_104,_zz_sbuf_wdat_4_105}}}};
  assign _zz_sbuf_wdat_4_10 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_11 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_12,_zz_sbuf_wdat_4_13}}}};
  assign _zz_sbuf_wdat_4_42 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_43 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_44,_zz_sbuf_wdat_4_45}}}};
  assign _zz_sbuf_wdat_4_74 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_75 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_76,_zz_sbuf_wdat_4_77}}}};
  assign _zz_sbuf_wdat_4_104 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_105 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_106,_zz_sbuf_wdat_4_107}}}};
  assign _zz_sbuf_wdat_4_12 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_13 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_14,_zz_sbuf_wdat_4_15}}}};
  assign _zz_sbuf_wdat_4_44 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_45 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_46,_zz_sbuf_wdat_4_47}}}};
  assign _zz_sbuf_wdat_4_76 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_77 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_78,_zz_sbuf_wdat_4_79}}}};
  assign _zz_sbuf_wdat_4_106 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_107 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_108,_zz_sbuf_wdat_4_109}}}};
  assign _zz_sbuf_wdat_4_14 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_15 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_16,_zz_sbuf_wdat_4_17}}}};
  assign _zz_sbuf_wdat_4_46 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_47 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_48,_zz_sbuf_wdat_4_49}}}};
  assign _zz_sbuf_wdat_4_78 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_79 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_80,_zz_sbuf_wdat_4_81}}}};
  assign _zz_sbuf_wdat_4_108 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_109 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_110,_zz_sbuf_wdat_4_111}}}};
  assign _zz_sbuf_wdat_4_16 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_17 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_18,_zz_sbuf_wdat_4_19}}}};
  assign _zz_sbuf_wdat_4_48 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_49 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_50,_zz_sbuf_wdat_4_51}}}};
  assign _zz_sbuf_wdat_4_80 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_81 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_82,_zz_sbuf_wdat_4_83}}}};
  assign _zz_sbuf_wdat_4_110 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_111 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_112,_zz_sbuf_wdat_4_113}}}};
  assign _zz_sbuf_wdat_4_18 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_19 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_20,_zz_sbuf_wdat_4_21}}}};
  assign _zz_sbuf_wdat_4_50 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_51 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_52,_zz_sbuf_wdat_4_53}}}};
  assign _zz_sbuf_wdat_4_82 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_83 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_84,_zz_sbuf_wdat_4_85}}}};
  assign _zz_sbuf_wdat_4_112 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_113 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_114,_zz_sbuf_wdat_4_115}}}};
  assign _zz_sbuf_wdat_4_20 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_21 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_22,_zz_sbuf_wdat_4_23}}}};
  assign _zz_sbuf_wdat_4_52 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_53 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_54,_zz_sbuf_wdat_4_55}}}};
  assign _zz_sbuf_wdat_4_84 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_85 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_86,_zz_sbuf_wdat_4_87}}}};
  assign _zz_sbuf_wdat_4_114 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_115 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_116,_zz_sbuf_wdat_4_117}}}};
  assign _zz_sbuf_wdat_4_22 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_23 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_24,_zz_sbuf_wdat_4_25}}}};
  assign _zz_sbuf_wdat_4_54 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_55 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_56,_zz_sbuf_wdat_4_57}}}};
  assign _zz_sbuf_wdat_4_86 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_87 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_88,_zz_sbuf_wdat_4_89}}}};
  assign _zz_sbuf_wdat_4_116 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_117 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_118,_zz_sbuf_wdat_4_119}}}};
  assign _zz_sbuf_wdat_4_24 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_25 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_26,_zz_sbuf_wdat_4_27}}}};
  assign _zz_sbuf_wdat_4_56 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_57 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_58,_zz_sbuf_wdat_4_59}}}};
  assign _zz_sbuf_wdat_4_88 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_89 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_90,_zz_sbuf_wdat_4_91}}}};
  assign _zz_sbuf_wdat_4_118 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_119 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_120,_zz_sbuf_wdat_4_121}}}};
  assign _zz_sbuf_wdat_4_26 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_27 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_28,_zz_sbuf_wdat_4_29}}}};
  assign _zz_sbuf_wdat_4_58 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_59 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_60,_zz_sbuf_wdat_4_61}}}};
  assign _zz_sbuf_wdat_4_90 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_91 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_92,_zz_sbuf_wdat_4_93}}}};
  assign _zz_sbuf_wdat_4_120 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_121 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_122,_zz_sbuf_wdat_4_123}}}};
  assign _zz_sbuf_wdat_4_28 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_29 = {dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_30,_zz_sbuf_wdat_4_31}}}}};
  assign _zz_sbuf_wdat_4_60 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_61 = {dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_62,_zz_sbuf_wdat_4_63}}}}};
  assign _zz_sbuf_wdat_4_92 = img2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_93 = {img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,img2sbuf_p0_wr_sel_4}}}};
  assign _zz_sbuf_wdat_4_122 = img2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_123 = {img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,img2sbuf_p1_wr_sel_4}}};
  assign _zz_sbuf_wdat_4_30 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_31 = dc2sbuf_p0_wr_sel_4;
  assign _zz_sbuf_wdat_4_62 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_4_63 = dc2sbuf_p1_wr_sel_4;
  assign _zz_sbuf_wdat_5 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_1 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_2,_zz_sbuf_wdat_5_3}}}};
  assign _zz_sbuf_wdat_5_32 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_33 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_34,_zz_sbuf_wdat_5_35}}}};
  assign _zz_sbuf_wdat_5_64 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_65 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_66,_zz_sbuf_wdat_5_67}}}};
  assign _zz_sbuf_wdat_5_94 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_95 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_96,_zz_sbuf_wdat_5_97}}}};
  assign _zz_sbuf_wdat_5_2 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_3 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_4,_zz_sbuf_wdat_5_5}}}};
  assign _zz_sbuf_wdat_5_34 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_35 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_36,_zz_sbuf_wdat_5_37}}}};
  assign _zz_sbuf_wdat_5_66 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_67 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_68,_zz_sbuf_wdat_5_69}}}};
  assign _zz_sbuf_wdat_5_96 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_97 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_98,_zz_sbuf_wdat_5_99}}}};
  assign _zz_sbuf_wdat_5_4 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_5 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_6,_zz_sbuf_wdat_5_7}}}};
  assign _zz_sbuf_wdat_5_36 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_37 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_38,_zz_sbuf_wdat_5_39}}}};
  assign _zz_sbuf_wdat_5_68 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_69 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_70,_zz_sbuf_wdat_5_71}}}};
  assign _zz_sbuf_wdat_5_98 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_99 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_100,_zz_sbuf_wdat_5_101}}}};
  assign _zz_sbuf_wdat_5_6 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_7 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_8,_zz_sbuf_wdat_5_9}}}};
  assign _zz_sbuf_wdat_5_38 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_39 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_40,_zz_sbuf_wdat_5_41}}}};
  assign _zz_sbuf_wdat_5_70 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_71 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_72,_zz_sbuf_wdat_5_73}}}};
  assign _zz_sbuf_wdat_5_100 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_101 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_102,_zz_sbuf_wdat_5_103}}}};
  assign _zz_sbuf_wdat_5_8 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_9 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_10,_zz_sbuf_wdat_5_11}}}};
  assign _zz_sbuf_wdat_5_40 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_41 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_42,_zz_sbuf_wdat_5_43}}}};
  assign _zz_sbuf_wdat_5_72 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_73 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_74,_zz_sbuf_wdat_5_75}}}};
  assign _zz_sbuf_wdat_5_102 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_103 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_104,_zz_sbuf_wdat_5_105}}}};
  assign _zz_sbuf_wdat_5_10 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_11 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_12,_zz_sbuf_wdat_5_13}}}};
  assign _zz_sbuf_wdat_5_42 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_43 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_44,_zz_sbuf_wdat_5_45}}}};
  assign _zz_sbuf_wdat_5_74 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_75 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_76,_zz_sbuf_wdat_5_77}}}};
  assign _zz_sbuf_wdat_5_104 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_105 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_106,_zz_sbuf_wdat_5_107}}}};
  assign _zz_sbuf_wdat_5_12 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_13 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_14,_zz_sbuf_wdat_5_15}}}};
  assign _zz_sbuf_wdat_5_44 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_45 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_46,_zz_sbuf_wdat_5_47}}}};
  assign _zz_sbuf_wdat_5_76 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_77 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_78,_zz_sbuf_wdat_5_79}}}};
  assign _zz_sbuf_wdat_5_106 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_107 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_108,_zz_sbuf_wdat_5_109}}}};
  assign _zz_sbuf_wdat_5_14 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_15 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_16,_zz_sbuf_wdat_5_17}}}};
  assign _zz_sbuf_wdat_5_46 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_47 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_48,_zz_sbuf_wdat_5_49}}}};
  assign _zz_sbuf_wdat_5_78 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_79 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_80,_zz_sbuf_wdat_5_81}}}};
  assign _zz_sbuf_wdat_5_108 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_109 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_110,_zz_sbuf_wdat_5_111}}}};
  assign _zz_sbuf_wdat_5_16 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_17 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_18,_zz_sbuf_wdat_5_19}}}};
  assign _zz_sbuf_wdat_5_48 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_49 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_50,_zz_sbuf_wdat_5_51}}}};
  assign _zz_sbuf_wdat_5_80 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_81 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_82,_zz_sbuf_wdat_5_83}}}};
  assign _zz_sbuf_wdat_5_110 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_111 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_112,_zz_sbuf_wdat_5_113}}}};
  assign _zz_sbuf_wdat_5_18 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_19 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_20,_zz_sbuf_wdat_5_21}}}};
  assign _zz_sbuf_wdat_5_50 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_51 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_52,_zz_sbuf_wdat_5_53}}}};
  assign _zz_sbuf_wdat_5_82 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_83 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_84,_zz_sbuf_wdat_5_85}}}};
  assign _zz_sbuf_wdat_5_112 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_113 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_114,_zz_sbuf_wdat_5_115}}}};
  assign _zz_sbuf_wdat_5_20 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_21 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_22,_zz_sbuf_wdat_5_23}}}};
  assign _zz_sbuf_wdat_5_52 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_53 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_54,_zz_sbuf_wdat_5_55}}}};
  assign _zz_sbuf_wdat_5_84 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_85 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_86,_zz_sbuf_wdat_5_87}}}};
  assign _zz_sbuf_wdat_5_114 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_115 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_116,_zz_sbuf_wdat_5_117}}}};
  assign _zz_sbuf_wdat_5_22 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_23 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_24,_zz_sbuf_wdat_5_25}}}};
  assign _zz_sbuf_wdat_5_54 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_55 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_56,_zz_sbuf_wdat_5_57}}}};
  assign _zz_sbuf_wdat_5_86 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_87 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_88,_zz_sbuf_wdat_5_89}}}};
  assign _zz_sbuf_wdat_5_116 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_117 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_118,_zz_sbuf_wdat_5_119}}}};
  assign _zz_sbuf_wdat_5_24 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_25 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_26,_zz_sbuf_wdat_5_27}}}};
  assign _zz_sbuf_wdat_5_56 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_57 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_58,_zz_sbuf_wdat_5_59}}}};
  assign _zz_sbuf_wdat_5_88 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_89 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_90,_zz_sbuf_wdat_5_91}}}};
  assign _zz_sbuf_wdat_5_118 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_119 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_120,_zz_sbuf_wdat_5_121}}}};
  assign _zz_sbuf_wdat_5_26 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_27 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_28,_zz_sbuf_wdat_5_29}}}};
  assign _zz_sbuf_wdat_5_58 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_59 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_60,_zz_sbuf_wdat_5_61}}}};
  assign _zz_sbuf_wdat_5_90 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_91 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_92,_zz_sbuf_wdat_5_93}}}};
  assign _zz_sbuf_wdat_5_120 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_121 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_122,_zz_sbuf_wdat_5_123}}}};
  assign _zz_sbuf_wdat_5_28 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_29 = {dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_30,_zz_sbuf_wdat_5_31}}}}};
  assign _zz_sbuf_wdat_5_60 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_61 = {dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_62,_zz_sbuf_wdat_5_63}}}}};
  assign _zz_sbuf_wdat_5_92 = img2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_93 = {img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,img2sbuf_p0_wr_sel_5}}}};
  assign _zz_sbuf_wdat_5_122 = img2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_123 = {img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,img2sbuf_p1_wr_sel_5}}};
  assign _zz_sbuf_wdat_5_30 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_31 = dc2sbuf_p0_wr_sel_5;
  assign _zz_sbuf_wdat_5_62 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_5_63 = dc2sbuf_p1_wr_sel_5;
  assign _zz_sbuf_wdat_6 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_1 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_2,_zz_sbuf_wdat_6_3}}}};
  assign _zz_sbuf_wdat_6_32 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_33 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_34,_zz_sbuf_wdat_6_35}}}};
  assign _zz_sbuf_wdat_6_64 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_65 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_66,_zz_sbuf_wdat_6_67}}}};
  assign _zz_sbuf_wdat_6_94 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_95 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_96,_zz_sbuf_wdat_6_97}}}};
  assign _zz_sbuf_wdat_6_2 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_3 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_4,_zz_sbuf_wdat_6_5}}}};
  assign _zz_sbuf_wdat_6_34 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_35 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_36,_zz_sbuf_wdat_6_37}}}};
  assign _zz_sbuf_wdat_6_66 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_67 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_68,_zz_sbuf_wdat_6_69}}}};
  assign _zz_sbuf_wdat_6_96 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_97 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_98,_zz_sbuf_wdat_6_99}}}};
  assign _zz_sbuf_wdat_6_4 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_5 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_6,_zz_sbuf_wdat_6_7}}}};
  assign _zz_sbuf_wdat_6_36 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_37 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_38,_zz_sbuf_wdat_6_39}}}};
  assign _zz_sbuf_wdat_6_68 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_69 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_70,_zz_sbuf_wdat_6_71}}}};
  assign _zz_sbuf_wdat_6_98 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_99 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_100,_zz_sbuf_wdat_6_101}}}};
  assign _zz_sbuf_wdat_6_6 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_7 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_8,_zz_sbuf_wdat_6_9}}}};
  assign _zz_sbuf_wdat_6_38 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_39 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_40,_zz_sbuf_wdat_6_41}}}};
  assign _zz_sbuf_wdat_6_70 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_71 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_72,_zz_sbuf_wdat_6_73}}}};
  assign _zz_sbuf_wdat_6_100 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_101 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_102,_zz_sbuf_wdat_6_103}}}};
  assign _zz_sbuf_wdat_6_8 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_9 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_10,_zz_sbuf_wdat_6_11}}}};
  assign _zz_sbuf_wdat_6_40 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_41 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_42,_zz_sbuf_wdat_6_43}}}};
  assign _zz_sbuf_wdat_6_72 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_73 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_74,_zz_sbuf_wdat_6_75}}}};
  assign _zz_sbuf_wdat_6_102 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_103 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_104,_zz_sbuf_wdat_6_105}}}};
  assign _zz_sbuf_wdat_6_10 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_11 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_12,_zz_sbuf_wdat_6_13}}}};
  assign _zz_sbuf_wdat_6_42 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_43 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_44,_zz_sbuf_wdat_6_45}}}};
  assign _zz_sbuf_wdat_6_74 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_75 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_76,_zz_sbuf_wdat_6_77}}}};
  assign _zz_sbuf_wdat_6_104 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_105 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_106,_zz_sbuf_wdat_6_107}}}};
  assign _zz_sbuf_wdat_6_12 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_13 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_14,_zz_sbuf_wdat_6_15}}}};
  assign _zz_sbuf_wdat_6_44 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_45 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_46,_zz_sbuf_wdat_6_47}}}};
  assign _zz_sbuf_wdat_6_76 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_77 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_78,_zz_sbuf_wdat_6_79}}}};
  assign _zz_sbuf_wdat_6_106 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_107 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_108,_zz_sbuf_wdat_6_109}}}};
  assign _zz_sbuf_wdat_6_14 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_15 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_16,_zz_sbuf_wdat_6_17}}}};
  assign _zz_sbuf_wdat_6_46 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_47 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_48,_zz_sbuf_wdat_6_49}}}};
  assign _zz_sbuf_wdat_6_78 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_79 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_80,_zz_sbuf_wdat_6_81}}}};
  assign _zz_sbuf_wdat_6_108 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_109 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_110,_zz_sbuf_wdat_6_111}}}};
  assign _zz_sbuf_wdat_6_16 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_17 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_18,_zz_sbuf_wdat_6_19}}}};
  assign _zz_sbuf_wdat_6_48 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_49 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_50,_zz_sbuf_wdat_6_51}}}};
  assign _zz_sbuf_wdat_6_80 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_81 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_82,_zz_sbuf_wdat_6_83}}}};
  assign _zz_sbuf_wdat_6_110 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_111 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_112,_zz_sbuf_wdat_6_113}}}};
  assign _zz_sbuf_wdat_6_18 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_19 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_20,_zz_sbuf_wdat_6_21}}}};
  assign _zz_sbuf_wdat_6_50 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_51 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_52,_zz_sbuf_wdat_6_53}}}};
  assign _zz_sbuf_wdat_6_82 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_83 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_84,_zz_sbuf_wdat_6_85}}}};
  assign _zz_sbuf_wdat_6_112 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_113 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_114,_zz_sbuf_wdat_6_115}}}};
  assign _zz_sbuf_wdat_6_20 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_21 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_22,_zz_sbuf_wdat_6_23}}}};
  assign _zz_sbuf_wdat_6_52 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_53 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_54,_zz_sbuf_wdat_6_55}}}};
  assign _zz_sbuf_wdat_6_84 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_85 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_86,_zz_sbuf_wdat_6_87}}}};
  assign _zz_sbuf_wdat_6_114 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_115 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_116,_zz_sbuf_wdat_6_117}}}};
  assign _zz_sbuf_wdat_6_22 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_23 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_24,_zz_sbuf_wdat_6_25}}}};
  assign _zz_sbuf_wdat_6_54 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_55 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_56,_zz_sbuf_wdat_6_57}}}};
  assign _zz_sbuf_wdat_6_86 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_87 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_88,_zz_sbuf_wdat_6_89}}}};
  assign _zz_sbuf_wdat_6_116 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_117 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_118,_zz_sbuf_wdat_6_119}}}};
  assign _zz_sbuf_wdat_6_24 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_25 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_26,_zz_sbuf_wdat_6_27}}}};
  assign _zz_sbuf_wdat_6_56 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_57 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_58,_zz_sbuf_wdat_6_59}}}};
  assign _zz_sbuf_wdat_6_88 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_89 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_90,_zz_sbuf_wdat_6_91}}}};
  assign _zz_sbuf_wdat_6_118 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_119 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_120,_zz_sbuf_wdat_6_121}}}};
  assign _zz_sbuf_wdat_6_26 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_27 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_28,_zz_sbuf_wdat_6_29}}}};
  assign _zz_sbuf_wdat_6_58 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_59 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_60,_zz_sbuf_wdat_6_61}}}};
  assign _zz_sbuf_wdat_6_90 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_91 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_92,_zz_sbuf_wdat_6_93}}}};
  assign _zz_sbuf_wdat_6_120 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_121 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_122,_zz_sbuf_wdat_6_123}}}};
  assign _zz_sbuf_wdat_6_28 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_29 = {dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_30,_zz_sbuf_wdat_6_31}}}}};
  assign _zz_sbuf_wdat_6_60 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_61 = {dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_62,_zz_sbuf_wdat_6_63}}}}};
  assign _zz_sbuf_wdat_6_92 = img2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_93 = {img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,img2sbuf_p0_wr_sel_6}}}};
  assign _zz_sbuf_wdat_6_122 = img2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_123 = {img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,img2sbuf_p1_wr_sel_6}}};
  assign _zz_sbuf_wdat_6_30 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_31 = dc2sbuf_p0_wr_sel_6;
  assign _zz_sbuf_wdat_6_62 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_6_63 = dc2sbuf_p1_wr_sel_6;
  assign _zz_sbuf_wdat_7 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_1 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_2,_zz_sbuf_wdat_7_3}}}};
  assign _zz_sbuf_wdat_7_32 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_33 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_34,_zz_sbuf_wdat_7_35}}}};
  assign _zz_sbuf_wdat_7_64 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_65 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_66,_zz_sbuf_wdat_7_67}}}};
  assign _zz_sbuf_wdat_7_94 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_95 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_96,_zz_sbuf_wdat_7_97}}}};
  assign _zz_sbuf_wdat_7_2 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_3 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_4,_zz_sbuf_wdat_7_5}}}};
  assign _zz_sbuf_wdat_7_34 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_35 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_36,_zz_sbuf_wdat_7_37}}}};
  assign _zz_sbuf_wdat_7_66 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_67 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_68,_zz_sbuf_wdat_7_69}}}};
  assign _zz_sbuf_wdat_7_96 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_97 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_98,_zz_sbuf_wdat_7_99}}}};
  assign _zz_sbuf_wdat_7_4 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_5 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_6,_zz_sbuf_wdat_7_7}}}};
  assign _zz_sbuf_wdat_7_36 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_37 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_38,_zz_sbuf_wdat_7_39}}}};
  assign _zz_sbuf_wdat_7_68 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_69 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_70,_zz_sbuf_wdat_7_71}}}};
  assign _zz_sbuf_wdat_7_98 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_99 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_100,_zz_sbuf_wdat_7_101}}}};
  assign _zz_sbuf_wdat_7_6 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_7 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_8,_zz_sbuf_wdat_7_9}}}};
  assign _zz_sbuf_wdat_7_38 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_39 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_40,_zz_sbuf_wdat_7_41}}}};
  assign _zz_sbuf_wdat_7_70 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_71 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_72,_zz_sbuf_wdat_7_73}}}};
  assign _zz_sbuf_wdat_7_100 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_101 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_102,_zz_sbuf_wdat_7_103}}}};
  assign _zz_sbuf_wdat_7_8 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_9 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_10,_zz_sbuf_wdat_7_11}}}};
  assign _zz_sbuf_wdat_7_40 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_41 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_42,_zz_sbuf_wdat_7_43}}}};
  assign _zz_sbuf_wdat_7_72 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_73 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_74,_zz_sbuf_wdat_7_75}}}};
  assign _zz_sbuf_wdat_7_102 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_103 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_104,_zz_sbuf_wdat_7_105}}}};
  assign _zz_sbuf_wdat_7_10 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_11 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_12,_zz_sbuf_wdat_7_13}}}};
  assign _zz_sbuf_wdat_7_42 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_43 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_44,_zz_sbuf_wdat_7_45}}}};
  assign _zz_sbuf_wdat_7_74 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_75 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_76,_zz_sbuf_wdat_7_77}}}};
  assign _zz_sbuf_wdat_7_104 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_105 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_106,_zz_sbuf_wdat_7_107}}}};
  assign _zz_sbuf_wdat_7_12 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_13 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_14,_zz_sbuf_wdat_7_15}}}};
  assign _zz_sbuf_wdat_7_44 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_45 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_46,_zz_sbuf_wdat_7_47}}}};
  assign _zz_sbuf_wdat_7_76 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_77 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_78,_zz_sbuf_wdat_7_79}}}};
  assign _zz_sbuf_wdat_7_106 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_107 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_108,_zz_sbuf_wdat_7_109}}}};
  assign _zz_sbuf_wdat_7_14 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_15 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_16,_zz_sbuf_wdat_7_17}}}};
  assign _zz_sbuf_wdat_7_46 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_47 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_48,_zz_sbuf_wdat_7_49}}}};
  assign _zz_sbuf_wdat_7_78 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_79 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_80,_zz_sbuf_wdat_7_81}}}};
  assign _zz_sbuf_wdat_7_108 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_109 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_110,_zz_sbuf_wdat_7_111}}}};
  assign _zz_sbuf_wdat_7_16 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_17 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_18,_zz_sbuf_wdat_7_19}}}};
  assign _zz_sbuf_wdat_7_48 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_49 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_50,_zz_sbuf_wdat_7_51}}}};
  assign _zz_sbuf_wdat_7_80 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_81 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_82,_zz_sbuf_wdat_7_83}}}};
  assign _zz_sbuf_wdat_7_110 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_111 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_112,_zz_sbuf_wdat_7_113}}}};
  assign _zz_sbuf_wdat_7_18 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_19 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_20,_zz_sbuf_wdat_7_21}}}};
  assign _zz_sbuf_wdat_7_50 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_51 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_52,_zz_sbuf_wdat_7_53}}}};
  assign _zz_sbuf_wdat_7_82 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_83 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_84,_zz_sbuf_wdat_7_85}}}};
  assign _zz_sbuf_wdat_7_112 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_113 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_114,_zz_sbuf_wdat_7_115}}}};
  assign _zz_sbuf_wdat_7_20 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_21 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_22,_zz_sbuf_wdat_7_23}}}};
  assign _zz_sbuf_wdat_7_52 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_53 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_54,_zz_sbuf_wdat_7_55}}}};
  assign _zz_sbuf_wdat_7_84 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_85 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_86,_zz_sbuf_wdat_7_87}}}};
  assign _zz_sbuf_wdat_7_114 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_115 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_116,_zz_sbuf_wdat_7_117}}}};
  assign _zz_sbuf_wdat_7_22 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_23 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_24,_zz_sbuf_wdat_7_25}}}};
  assign _zz_sbuf_wdat_7_54 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_55 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_56,_zz_sbuf_wdat_7_57}}}};
  assign _zz_sbuf_wdat_7_86 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_87 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_88,_zz_sbuf_wdat_7_89}}}};
  assign _zz_sbuf_wdat_7_116 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_117 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_118,_zz_sbuf_wdat_7_119}}}};
  assign _zz_sbuf_wdat_7_24 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_25 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_26,_zz_sbuf_wdat_7_27}}}};
  assign _zz_sbuf_wdat_7_56 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_57 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_58,_zz_sbuf_wdat_7_59}}}};
  assign _zz_sbuf_wdat_7_88 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_89 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_90,_zz_sbuf_wdat_7_91}}}};
  assign _zz_sbuf_wdat_7_118 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_119 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_120,_zz_sbuf_wdat_7_121}}}};
  assign _zz_sbuf_wdat_7_26 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_27 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_28,_zz_sbuf_wdat_7_29}}}};
  assign _zz_sbuf_wdat_7_58 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_59 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_60,_zz_sbuf_wdat_7_61}}}};
  assign _zz_sbuf_wdat_7_90 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_91 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_92,_zz_sbuf_wdat_7_93}}}};
  assign _zz_sbuf_wdat_7_120 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_121 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_122,_zz_sbuf_wdat_7_123}}}};
  assign _zz_sbuf_wdat_7_28 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_29 = {dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_30,_zz_sbuf_wdat_7_31}}}}};
  assign _zz_sbuf_wdat_7_60 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_61 = {dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_62,_zz_sbuf_wdat_7_63}}}}};
  assign _zz_sbuf_wdat_7_92 = img2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_93 = {img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,img2sbuf_p0_wr_sel_7}}}};
  assign _zz_sbuf_wdat_7_122 = img2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_123 = {img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,img2sbuf_p1_wr_sel_7}}};
  assign _zz_sbuf_wdat_7_30 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_31 = dc2sbuf_p0_wr_sel_7;
  assign _zz_sbuf_wdat_7_62 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_7_63 = dc2sbuf_p1_wr_sel_7;
  assign _zz_sbuf_wdat_8 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_1 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_2,_zz_sbuf_wdat_8_3}}}};
  assign _zz_sbuf_wdat_8_32 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_33 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_34,_zz_sbuf_wdat_8_35}}}};
  assign _zz_sbuf_wdat_8_64 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_65 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_66,_zz_sbuf_wdat_8_67}}}};
  assign _zz_sbuf_wdat_8_94 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_95 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_96,_zz_sbuf_wdat_8_97}}}};
  assign _zz_sbuf_wdat_8_2 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_3 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_4,_zz_sbuf_wdat_8_5}}}};
  assign _zz_sbuf_wdat_8_34 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_35 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_36,_zz_sbuf_wdat_8_37}}}};
  assign _zz_sbuf_wdat_8_66 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_67 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_68,_zz_sbuf_wdat_8_69}}}};
  assign _zz_sbuf_wdat_8_96 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_97 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_98,_zz_sbuf_wdat_8_99}}}};
  assign _zz_sbuf_wdat_8_4 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_5 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_6,_zz_sbuf_wdat_8_7}}}};
  assign _zz_sbuf_wdat_8_36 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_37 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_38,_zz_sbuf_wdat_8_39}}}};
  assign _zz_sbuf_wdat_8_68 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_69 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_70,_zz_sbuf_wdat_8_71}}}};
  assign _zz_sbuf_wdat_8_98 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_99 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_100,_zz_sbuf_wdat_8_101}}}};
  assign _zz_sbuf_wdat_8_6 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_7 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_8,_zz_sbuf_wdat_8_9}}}};
  assign _zz_sbuf_wdat_8_38 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_39 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_40,_zz_sbuf_wdat_8_41}}}};
  assign _zz_sbuf_wdat_8_70 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_71 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_72,_zz_sbuf_wdat_8_73}}}};
  assign _zz_sbuf_wdat_8_100 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_101 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_102,_zz_sbuf_wdat_8_103}}}};
  assign _zz_sbuf_wdat_8_8 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_9 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_10,_zz_sbuf_wdat_8_11}}}};
  assign _zz_sbuf_wdat_8_40 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_41 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_42,_zz_sbuf_wdat_8_43}}}};
  assign _zz_sbuf_wdat_8_72 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_73 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_74,_zz_sbuf_wdat_8_75}}}};
  assign _zz_sbuf_wdat_8_102 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_103 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_104,_zz_sbuf_wdat_8_105}}}};
  assign _zz_sbuf_wdat_8_10 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_11 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_12,_zz_sbuf_wdat_8_13}}}};
  assign _zz_sbuf_wdat_8_42 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_43 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_44,_zz_sbuf_wdat_8_45}}}};
  assign _zz_sbuf_wdat_8_74 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_75 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_76,_zz_sbuf_wdat_8_77}}}};
  assign _zz_sbuf_wdat_8_104 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_105 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_106,_zz_sbuf_wdat_8_107}}}};
  assign _zz_sbuf_wdat_8_12 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_13 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_14,_zz_sbuf_wdat_8_15}}}};
  assign _zz_sbuf_wdat_8_44 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_45 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_46,_zz_sbuf_wdat_8_47}}}};
  assign _zz_sbuf_wdat_8_76 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_77 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_78,_zz_sbuf_wdat_8_79}}}};
  assign _zz_sbuf_wdat_8_106 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_107 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_108,_zz_sbuf_wdat_8_109}}}};
  assign _zz_sbuf_wdat_8_14 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_15 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_16,_zz_sbuf_wdat_8_17}}}};
  assign _zz_sbuf_wdat_8_46 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_47 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_48,_zz_sbuf_wdat_8_49}}}};
  assign _zz_sbuf_wdat_8_78 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_79 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_80,_zz_sbuf_wdat_8_81}}}};
  assign _zz_sbuf_wdat_8_108 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_109 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_110,_zz_sbuf_wdat_8_111}}}};
  assign _zz_sbuf_wdat_8_16 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_17 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_18,_zz_sbuf_wdat_8_19}}}};
  assign _zz_sbuf_wdat_8_48 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_49 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_50,_zz_sbuf_wdat_8_51}}}};
  assign _zz_sbuf_wdat_8_80 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_81 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_82,_zz_sbuf_wdat_8_83}}}};
  assign _zz_sbuf_wdat_8_110 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_111 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_112,_zz_sbuf_wdat_8_113}}}};
  assign _zz_sbuf_wdat_8_18 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_19 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_20,_zz_sbuf_wdat_8_21}}}};
  assign _zz_sbuf_wdat_8_50 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_51 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_52,_zz_sbuf_wdat_8_53}}}};
  assign _zz_sbuf_wdat_8_82 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_83 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_84,_zz_sbuf_wdat_8_85}}}};
  assign _zz_sbuf_wdat_8_112 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_113 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_114,_zz_sbuf_wdat_8_115}}}};
  assign _zz_sbuf_wdat_8_20 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_21 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_22,_zz_sbuf_wdat_8_23}}}};
  assign _zz_sbuf_wdat_8_52 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_53 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_54,_zz_sbuf_wdat_8_55}}}};
  assign _zz_sbuf_wdat_8_84 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_85 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_86,_zz_sbuf_wdat_8_87}}}};
  assign _zz_sbuf_wdat_8_114 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_115 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_116,_zz_sbuf_wdat_8_117}}}};
  assign _zz_sbuf_wdat_8_22 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_23 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_24,_zz_sbuf_wdat_8_25}}}};
  assign _zz_sbuf_wdat_8_54 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_55 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_56,_zz_sbuf_wdat_8_57}}}};
  assign _zz_sbuf_wdat_8_86 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_87 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_88,_zz_sbuf_wdat_8_89}}}};
  assign _zz_sbuf_wdat_8_116 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_117 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_118,_zz_sbuf_wdat_8_119}}}};
  assign _zz_sbuf_wdat_8_24 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_25 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_26,_zz_sbuf_wdat_8_27}}}};
  assign _zz_sbuf_wdat_8_56 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_57 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_58,_zz_sbuf_wdat_8_59}}}};
  assign _zz_sbuf_wdat_8_88 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_89 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_90,_zz_sbuf_wdat_8_91}}}};
  assign _zz_sbuf_wdat_8_118 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_119 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_120,_zz_sbuf_wdat_8_121}}}};
  assign _zz_sbuf_wdat_8_26 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_27 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_28,_zz_sbuf_wdat_8_29}}}};
  assign _zz_sbuf_wdat_8_58 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_59 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_60,_zz_sbuf_wdat_8_61}}}};
  assign _zz_sbuf_wdat_8_90 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_91 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_92,_zz_sbuf_wdat_8_93}}}};
  assign _zz_sbuf_wdat_8_120 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_121 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_122,_zz_sbuf_wdat_8_123}}}};
  assign _zz_sbuf_wdat_8_28 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_29 = {dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_30,_zz_sbuf_wdat_8_31}}}}};
  assign _zz_sbuf_wdat_8_60 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_61 = {dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_62,_zz_sbuf_wdat_8_63}}}}};
  assign _zz_sbuf_wdat_8_92 = img2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_93 = {img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,img2sbuf_p0_wr_sel_8}}}};
  assign _zz_sbuf_wdat_8_122 = img2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_123 = {img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,img2sbuf_p1_wr_sel_8}}};
  assign _zz_sbuf_wdat_8_30 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_31 = dc2sbuf_p0_wr_sel_8;
  assign _zz_sbuf_wdat_8_62 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_8_63 = dc2sbuf_p1_wr_sel_8;
  assign _zz_sbuf_wdat_9 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_1 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_2,_zz_sbuf_wdat_9_3}}}};
  assign _zz_sbuf_wdat_9_32 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_33 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_34,_zz_sbuf_wdat_9_35}}}};
  assign _zz_sbuf_wdat_9_64 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_65 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_66,_zz_sbuf_wdat_9_67}}}};
  assign _zz_sbuf_wdat_9_94 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_95 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_96,_zz_sbuf_wdat_9_97}}}};
  assign _zz_sbuf_wdat_9_2 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_3 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_4,_zz_sbuf_wdat_9_5}}}};
  assign _zz_sbuf_wdat_9_34 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_35 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_36,_zz_sbuf_wdat_9_37}}}};
  assign _zz_sbuf_wdat_9_66 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_67 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_68,_zz_sbuf_wdat_9_69}}}};
  assign _zz_sbuf_wdat_9_96 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_97 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_98,_zz_sbuf_wdat_9_99}}}};
  assign _zz_sbuf_wdat_9_4 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_5 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_6,_zz_sbuf_wdat_9_7}}}};
  assign _zz_sbuf_wdat_9_36 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_37 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_38,_zz_sbuf_wdat_9_39}}}};
  assign _zz_sbuf_wdat_9_68 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_69 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_70,_zz_sbuf_wdat_9_71}}}};
  assign _zz_sbuf_wdat_9_98 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_99 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_100,_zz_sbuf_wdat_9_101}}}};
  assign _zz_sbuf_wdat_9_6 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_7 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_8,_zz_sbuf_wdat_9_9}}}};
  assign _zz_sbuf_wdat_9_38 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_39 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_40,_zz_sbuf_wdat_9_41}}}};
  assign _zz_sbuf_wdat_9_70 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_71 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_72,_zz_sbuf_wdat_9_73}}}};
  assign _zz_sbuf_wdat_9_100 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_101 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_102,_zz_sbuf_wdat_9_103}}}};
  assign _zz_sbuf_wdat_9_8 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_9 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_10,_zz_sbuf_wdat_9_11}}}};
  assign _zz_sbuf_wdat_9_40 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_41 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_42,_zz_sbuf_wdat_9_43}}}};
  assign _zz_sbuf_wdat_9_72 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_73 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_74,_zz_sbuf_wdat_9_75}}}};
  assign _zz_sbuf_wdat_9_102 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_103 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_104,_zz_sbuf_wdat_9_105}}}};
  assign _zz_sbuf_wdat_9_10 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_11 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_12,_zz_sbuf_wdat_9_13}}}};
  assign _zz_sbuf_wdat_9_42 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_43 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_44,_zz_sbuf_wdat_9_45}}}};
  assign _zz_sbuf_wdat_9_74 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_75 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_76,_zz_sbuf_wdat_9_77}}}};
  assign _zz_sbuf_wdat_9_104 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_105 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_106,_zz_sbuf_wdat_9_107}}}};
  assign _zz_sbuf_wdat_9_12 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_13 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_14,_zz_sbuf_wdat_9_15}}}};
  assign _zz_sbuf_wdat_9_44 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_45 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_46,_zz_sbuf_wdat_9_47}}}};
  assign _zz_sbuf_wdat_9_76 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_77 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_78,_zz_sbuf_wdat_9_79}}}};
  assign _zz_sbuf_wdat_9_106 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_107 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_108,_zz_sbuf_wdat_9_109}}}};
  assign _zz_sbuf_wdat_9_14 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_15 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_16,_zz_sbuf_wdat_9_17}}}};
  assign _zz_sbuf_wdat_9_46 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_47 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_48,_zz_sbuf_wdat_9_49}}}};
  assign _zz_sbuf_wdat_9_78 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_79 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_80,_zz_sbuf_wdat_9_81}}}};
  assign _zz_sbuf_wdat_9_108 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_109 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_110,_zz_sbuf_wdat_9_111}}}};
  assign _zz_sbuf_wdat_9_16 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_17 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_18,_zz_sbuf_wdat_9_19}}}};
  assign _zz_sbuf_wdat_9_48 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_49 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_50,_zz_sbuf_wdat_9_51}}}};
  assign _zz_sbuf_wdat_9_80 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_81 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_82,_zz_sbuf_wdat_9_83}}}};
  assign _zz_sbuf_wdat_9_110 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_111 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_112,_zz_sbuf_wdat_9_113}}}};
  assign _zz_sbuf_wdat_9_18 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_19 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_20,_zz_sbuf_wdat_9_21}}}};
  assign _zz_sbuf_wdat_9_50 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_51 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_52,_zz_sbuf_wdat_9_53}}}};
  assign _zz_sbuf_wdat_9_82 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_83 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_84,_zz_sbuf_wdat_9_85}}}};
  assign _zz_sbuf_wdat_9_112 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_113 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_114,_zz_sbuf_wdat_9_115}}}};
  assign _zz_sbuf_wdat_9_20 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_21 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_22,_zz_sbuf_wdat_9_23}}}};
  assign _zz_sbuf_wdat_9_52 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_53 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_54,_zz_sbuf_wdat_9_55}}}};
  assign _zz_sbuf_wdat_9_84 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_85 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_86,_zz_sbuf_wdat_9_87}}}};
  assign _zz_sbuf_wdat_9_114 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_115 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_116,_zz_sbuf_wdat_9_117}}}};
  assign _zz_sbuf_wdat_9_22 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_23 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_24,_zz_sbuf_wdat_9_25}}}};
  assign _zz_sbuf_wdat_9_54 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_55 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_56,_zz_sbuf_wdat_9_57}}}};
  assign _zz_sbuf_wdat_9_86 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_87 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_88,_zz_sbuf_wdat_9_89}}}};
  assign _zz_sbuf_wdat_9_116 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_117 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_118,_zz_sbuf_wdat_9_119}}}};
  assign _zz_sbuf_wdat_9_24 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_25 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_26,_zz_sbuf_wdat_9_27}}}};
  assign _zz_sbuf_wdat_9_56 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_57 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_58,_zz_sbuf_wdat_9_59}}}};
  assign _zz_sbuf_wdat_9_88 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_89 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_90,_zz_sbuf_wdat_9_91}}}};
  assign _zz_sbuf_wdat_9_118 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_119 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_120,_zz_sbuf_wdat_9_121}}}};
  assign _zz_sbuf_wdat_9_26 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_27 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_28,_zz_sbuf_wdat_9_29}}}};
  assign _zz_sbuf_wdat_9_58 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_59 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_60,_zz_sbuf_wdat_9_61}}}};
  assign _zz_sbuf_wdat_9_90 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_91 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_92,_zz_sbuf_wdat_9_93}}}};
  assign _zz_sbuf_wdat_9_120 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_121 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_122,_zz_sbuf_wdat_9_123}}}};
  assign _zz_sbuf_wdat_9_28 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_29 = {dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_30,_zz_sbuf_wdat_9_31}}}}};
  assign _zz_sbuf_wdat_9_60 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_61 = {dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_62,_zz_sbuf_wdat_9_63}}}}};
  assign _zz_sbuf_wdat_9_92 = img2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_93 = {img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,img2sbuf_p0_wr_sel_9}}}};
  assign _zz_sbuf_wdat_9_122 = img2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_123 = {img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,img2sbuf_p1_wr_sel_9}}};
  assign _zz_sbuf_wdat_9_30 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_31 = dc2sbuf_p0_wr_sel_9;
  assign _zz_sbuf_wdat_9_62 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_9_63 = dc2sbuf_p1_wr_sel_9;
  assign _zz_sbuf_wdat_10 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_1 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_2,_zz_sbuf_wdat_10_3}}}};
  assign _zz_sbuf_wdat_10_32 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_33 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_34,_zz_sbuf_wdat_10_35}}}};
  assign _zz_sbuf_wdat_10_64 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_65 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_66,_zz_sbuf_wdat_10_67}}}};
  assign _zz_sbuf_wdat_10_94 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_95 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_96,_zz_sbuf_wdat_10_97}}}};
  assign _zz_sbuf_wdat_10_2 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_3 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_4,_zz_sbuf_wdat_10_5}}}};
  assign _zz_sbuf_wdat_10_34 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_35 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_36,_zz_sbuf_wdat_10_37}}}};
  assign _zz_sbuf_wdat_10_66 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_67 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_68,_zz_sbuf_wdat_10_69}}}};
  assign _zz_sbuf_wdat_10_96 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_97 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_98,_zz_sbuf_wdat_10_99}}}};
  assign _zz_sbuf_wdat_10_4 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_5 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_6,_zz_sbuf_wdat_10_7}}}};
  assign _zz_sbuf_wdat_10_36 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_37 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_38,_zz_sbuf_wdat_10_39}}}};
  assign _zz_sbuf_wdat_10_68 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_69 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_70,_zz_sbuf_wdat_10_71}}}};
  assign _zz_sbuf_wdat_10_98 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_99 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_100,_zz_sbuf_wdat_10_101}}}};
  assign _zz_sbuf_wdat_10_6 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_7 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_8,_zz_sbuf_wdat_10_9}}}};
  assign _zz_sbuf_wdat_10_38 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_39 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_40,_zz_sbuf_wdat_10_41}}}};
  assign _zz_sbuf_wdat_10_70 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_71 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_72,_zz_sbuf_wdat_10_73}}}};
  assign _zz_sbuf_wdat_10_100 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_101 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_102,_zz_sbuf_wdat_10_103}}}};
  assign _zz_sbuf_wdat_10_8 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_9 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_10,_zz_sbuf_wdat_10_11}}}};
  assign _zz_sbuf_wdat_10_40 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_41 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_42,_zz_sbuf_wdat_10_43}}}};
  assign _zz_sbuf_wdat_10_72 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_73 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_74,_zz_sbuf_wdat_10_75}}}};
  assign _zz_sbuf_wdat_10_102 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_103 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_104,_zz_sbuf_wdat_10_105}}}};
  assign _zz_sbuf_wdat_10_10 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_11 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_12,_zz_sbuf_wdat_10_13}}}};
  assign _zz_sbuf_wdat_10_42 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_43 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_44,_zz_sbuf_wdat_10_45}}}};
  assign _zz_sbuf_wdat_10_74 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_75 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_76,_zz_sbuf_wdat_10_77}}}};
  assign _zz_sbuf_wdat_10_104 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_105 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_106,_zz_sbuf_wdat_10_107}}}};
  assign _zz_sbuf_wdat_10_12 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_13 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_14,_zz_sbuf_wdat_10_15}}}};
  assign _zz_sbuf_wdat_10_44 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_45 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_46,_zz_sbuf_wdat_10_47}}}};
  assign _zz_sbuf_wdat_10_76 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_77 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_78,_zz_sbuf_wdat_10_79}}}};
  assign _zz_sbuf_wdat_10_106 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_107 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_108,_zz_sbuf_wdat_10_109}}}};
  assign _zz_sbuf_wdat_10_14 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_15 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_16,_zz_sbuf_wdat_10_17}}}};
  assign _zz_sbuf_wdat_10_46 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_47 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_48,_zz_sbuf_wdat_10_49}}}};
  assign _zz_sbuf_wdat_10_78 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_79 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_80,_zz_sbuf_wdat_10_81}}}};
  assign _zz_sbuf_wdat_10_108 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_109 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_110,_zz_sbuf_wdat_10_111}}}};
  assign _zz_sbuf_wdat_10_16 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_17 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_18,_zz_sbuf_wdat_10_19}}}};
  assign _zz_sbuf_wdat_10_48 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_49 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_50,_zz_sbuf_wdat_10_51}}}};
  assign _zz_sbuf_wdat_10_80 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_81 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_82,_zz_sbuf_wdat_10_83}}}};
  assign _zz_sbuf_wdat_10_110 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_111 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_112,_zz_sbuf_wdat_10_113}}}};
  assign _zz_sbuf_wdat_10_18 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_19 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_20,_zz_sbuf_wdat_10_21}}}};
  assign _zz_sbuf_wdat_10_50 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_51 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_52,_zz_sbuf_wdat_10_53}}}};
  assign _zz_sbuf_wdat_10_82 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_83 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_84,_zz_sbuf_wdat_10_85}}}};
  assign _zz_sbuf_wdat_10_112 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_113 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_114,_zz_sbuf_wdat_10_115}}}};
  assign _zz_sbuf_wdat_10_20 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_21 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_22,_zz_sbuf_wdat_10_23}}}};
  assign _zz_sbuf_wdat_10_52 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_53 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_54,_zz_sbuf_wdat_10_55}}}};
  assign _zz_sbuf_wdat_10_84 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_85 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_86,_zz_sbuf_wdat_10_87}}}};
  assign _zz_sbuf_wdat_10_114 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_115 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_116,_zz_sbuf_wdat_10_117}}}};
  assign _zz_sbuf_wdat_10_22 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_23 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_24,_zz_sbuf_wdat_10_25}}}};
  assign _zz_sbuf_wdat_10_54 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_55 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_56,_zz_sbuf_wdat_10_57}}}};
  assign _zz_sbuf_wdat_10_86 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_87 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_88,_zz_sbuf_wdat_10_89}}}};
  assign _zz_sbuf_wdat_10_116 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_117 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_118,_zz_sbuf_wdat_10_119}}}};
  assign _zz_sbuf_wdat_10_24 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_25 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_26,_zz_sbuf_wdat_10_27}}}};
  assign _zz_sbuf_wdat_10_56 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_57 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_58,_zz_sbuf_wdat_10_59}}}};
  assign _zz_sbuf_wdat_10_88 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_89 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_90,_zz_sbuf_wdat_10_91}}}};
  assign _zz_sbuf_wdat_10_118 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_119 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_120,_zz_sbuf_wdat_10_121}}}};
  assign _zz_sbuf_wdat_10_26 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_27 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_28,_zz_sbuf_wdat_10_29}}}};
  assign _zz_sbuf_wdat_10_58 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_59 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_60,_zz_sbuf_wdat_10_61}}}};
  assign _zz_sbuf_wdat_10_90 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_91 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_92,_zz_sbuf_wdat_10_93}}}};
  assign _zz_sbuf_wdat_10_120 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_121 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_122,_zz_sbuf_wdat_10_123}}}};
  assign _zz_sbuf_wdat_10_28 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_29 = {dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_30,_zz_sbuf_wdat_10_31}}}}};
  assign _zz_sbuf_wdat_10_60 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_61 = {dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_62,_zz_sbuf_wdat_10_63}}}}};
  assign _zz_sbuf_wdat_10_92 = img2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_93 = {img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,img2sbuf_p0_wr_sel_10}}}};
  assign _zz_sbuf_wdat_10_122 = img2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_123 = {img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,img2sbuf_p1_wr_sel_10}}};
  assign _zz_sbuf_wdat_10_30 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_31 = dc2sbuf_p0_wr_sel_10;
  assign _zz_sbuf_wdat_10_62 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_10_63 = dc2sbuf_p1_wr_sel_10;
  assign _zz_sbuf_wdat_11 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_1 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_2,_zz_sbuf_wdat_11_3}}}};
  assign _zz_sbuf_wdat_11_32 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_33 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_34,_zz_sbuf_wdat_11_35}}}};
  assign _zz_sbuf_wdat_11_64 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_65 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_66,_zz_sbuf_wdat_11_67}}}};
  assign _zz_sbuf_wdat_11_94 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_95 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_96,_zz_sbuf_wdat_11_97}}}};
  assign _zz_sbuf_wdat_11_2 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_3 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_4,_zz_sbuf_wdat_11_5}}}};
  assign _zz_sbuf_wdat_11_34 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_35 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_36,_zz_sbuf_wdat_11_37}}}};
  assign _zz_sbuf_wdat_11_66 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_67 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_68,_zz_sbuf_wdat_11_69}}}};
  assign _zz_sbuf_wdat_11_96 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_97 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_98,_zz_sbuf_wdat_11_99}}}};
  assign _zz_sbuf_wdat_11_4 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_5 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_6,_zz_sbuf_wdat_11_7}}}};
  assign _zz_sbuf_wdat_11_36 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_37 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_38,_zz_sbuf_wdat_11_39}}}};
  assign _zz_sbuf_wdat_11_68 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_69 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_70,_zz_sbuf_wdat_11_71}}}};
  assign _zz_sbuf_wdat_11_98 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_99 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_100,_zz_sbuf_wdat_11_101}}}};
  assign _zz_sbuf_wdat_11_6 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_7 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_8,_zz_sbuf_wdat_11_9}}}};
  assign _zz_sbuf_wdat_11_38 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_39 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_40,_zz_sbuf_wdat_11_41}}}};
  assign _zz_sbuf_wdat_11_70 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_71 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_72,_zz_sbuf_wdat_11_73}}}};
  assign _zz_sbuf_wdat_11_100 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_101 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_102,_zz_sbuf_wdat_11_103}}}};
  assign _zz_sbuf_wdat_11_8 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_9 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_10,_zz_sbuf_wdat_11_11}}}};
  assign _zz_sbuf_wdat_11_40 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_41 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_42,_zz_sbuf_wdat_11_43}}}};
  assign _zz_sbuf_wdat_11_72 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_73 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_74,_zz_sbuf_wdat_11_75}}}};
  assign _zz_sbuf_wdat_11_102 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_103 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_104,_zz_sbuf_wdat_11_105}}}};
  assign _zz_sbuf_wdat_11_10 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_11 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_12,_zz_sbuf_wdat_11_13}}}};
  assign _zz_sbuf_wdat_11_42 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_43 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_44,_zz_sbuf_wdat_11_45}}}};
  assign _zz_sbuf_wdat_11_74 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_75 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_76,_zz_sbuf_wdat_11_77}}}};
  assign _zz_sbuf_wdat_11_104 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_105 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_106,_zz_sbuf_wdat_11_107}}}};
  assign _zz_sbuf_wdat_11_12 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_13 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_14,_zz_sbuf_wdat_11_15}}}};
  assign _zz_sbuf_wdat_11_44 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_45 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_46,_zz_sbuf_wdat_11_47}}}};
  assign _zz_sbuf_wdat_11_76 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_77 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_78,_zz_sbuf_wdat_11_79}}}};
  assign _zz_sbuf_wdat_11_106 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_107 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_108,_zz_sbuf_wdat_11_109}}}};
  assign _zz_sbuf_wdat_11_14 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_15 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_16,_zz_sbuf_wdat_11_17}}}};
  assign _zz_sbuf_wdat_11_46 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_47 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_48,_zz_sbuf_wdat_11_49}}}};
  assign _zz_sbuf_wdat_11_78 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_79 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_80,_zz_sbuf_wdat_11_81}}}};
  assign _zz_sbuf_wdat_11_108 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_109 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_110,_zz_sbuf_wdat_11_111}}}};
  assign _zz_sbuf_wdat_11_16 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_17 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_18,_zz_sbuf_wdat_11_19}}}};
  assign _zz_sbuf_wdat_11_48 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_49 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_50,_zz_sbuf_wdat_11_51}}}};
  assign _zz_sbuf_wdat_11_80 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_81 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_82,_zz_sbuf_wdat_11_83}}}};
  assign _zz_sbuf_wdat_11_110 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_111 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_112,_zz_sbuf_wdat_11_113}}}};
  assign _zz_sbuf_wdat_11_18 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_19 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_20,_zz_sbuf_wdat_11_21}}}};
  assign _zz_sbuf_wdat_11_50 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_51 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_52,_zz_sbuf_wdat_11_53}}}};
  assign _zz_sbuf_wdat_11_82 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_83 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_84,_zz_sbuf_wdat_11_85}}}};
  assign _zz_sbuf_wdat_11_112 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_113 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_114,_zz_sbuf_wdat_11_115}}}};
  assign _zz_sbuf_wdat_11_20 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_21 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_22,_zz_sbuf_wdat_11_23}}}};
  assign _zz_sbuf_wdat_11_52 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_53 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_54,_zz_sbuf_wdat_11_55}}}};
  assign _zz_sbuf_wdat_11_84 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_85 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_86,_zz_sbuf_wdat_11_87}}}};
  assign _zz_sbuf_wdat_11_114 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_115 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_116,_zz_sbuf_wdat_11_117}}}};
  assign _zz_sbuf_wdat_11_22 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_23 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_24,_zz_sbuf_wdat_11_25}}}};
  assign _zz_sbuf_wdat_11_54 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_55 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_56,_zz_sbuf_wdat_11_57}}}};
  assign _zz_sbuf_wdat_11_86 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_87 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_88,_zz_sbuf_wdat_11_89}}}};
  assign _zz_sbuf_wdat_11_116 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_117 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_118,_zz_sbuf_wdat_11_119}}}};
  assign _zz_sbuf_wdat_11_24 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_25 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_26,_zz_sbuf_wdat_11_27}}}};
  assign _zz_sbuf_wdat_11_56 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_57 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_58,_zz_sbuf_wdat_11_59}}}};
  assign _zz_sbuf_wdat_11_88 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_89 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_90,_zz_sbuf_wdat_11_91}}}};
  assign _zz_sbuf_wdat_11_118 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_119 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_120,_zz_sbuf_wdat_11_121}}}};
  assign _zz_sbuf_wdat_11_26 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_27 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_28,_zz_sbuf_wdat_11_29}}}};
  assign _zz_sbuf_wdat_11_58 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_59 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_60,_zz_sbuf_wdat_11_61}}}};
  assign _zz_sbuf_wdat_11_90 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_91 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_92,_zz_sbuf_wdat_11_93}}}};
  assign _zz_sbuf_wdat_11_120 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_121 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_122,_zz_sbuf_wdat_11_123}}}};
  assign _zz_sbuf_wdat_11_28 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_29 = {dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_30,_zz_sbuf_wdat_11_31}}}}};
  assign _zz_sbuf_wdat_11_60 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_61 = {dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_62,_zz_sbuf_wdat_11_63}}}}};
  assign _zz_sbuf_wdat_11_92 = img2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_93 = {img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,img2sbuf_p0_wr_sel_11}}}};
  assign _zz_sbuf_wdat_11_122 = img2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_123 = {img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,img2sbuf_p1_wr_sel_11}}};
  assign _zz_sbuf_wdat_11_30 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_31 = dc2sbuf_p0_wr_sel_11;
  assign _zz_sbuf_wdat_11_62 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_11_63 = dc2sbuf_p1_wr_sel_11;
  assign _zz_sbuf_wdat_12 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_1 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_2,_zz_sbuf_wdat_12_3}}}};
  assign _zz_sbuf_wdat_12_32 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_33 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_34,_zz_sbuf_wdat_12_35}}}};
  assign _zz_sbuf_wdat_12_64 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_65 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_66,_zz_sbuf_wdat_12_67}}}};
  assign _zz_sbuf_wdat_12_94 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_95 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_96,_zz_sbuf_wdat_12_97}}}};
  assign _zz_sbuf_wdat_12_2 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_3 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_4,_zz_sbuf_wdat_12_5}}}};
  assign _zz_sbuf_wdat_12_34 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_35 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_36,_zz_sbuf_wdat_12_37}}}};
  assign _zz_sbuf_wdat_12_66 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_67 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_68,_zz_sbuf_wdat_12_69}}}};
  assign _zz_sbuf_wdat_12_96 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_97 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_98,_zz_sbuf_wdat_12_99}}}};
  assign _zz_sbuf_wdat_12_4 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_5 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_6,_zz_sbuf_wdat_12_7}}}};
  assign _zz_sbuf_wdat_12_36 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_37 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_38,_zz_sbuf_wdat_12_39}}}};
  assign _zz_sbuf_wdat_12_68 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_69 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_70,_zz_sbuf_wdat_12_71}}}};
  assign _zz_sbuf_wdat_12_98 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_99 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_100,_zz_sbuf_wdat_12_101}}}};
  assign _zz_sbuf_wdat_12_6 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_7 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_8,_zz_sbuf_wdat_12_9}}}};
  assign _zz_sbuf_wdat_12_38 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_39 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_40,_zz_sbuf_wdat_12_41}}}};
  assign _zz_sbuf_wdat_12_70 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_71 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_72,_zz_sbuf_wdat_12_73}}}};
  assign _zz_sbuf_wdat_12_100 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_101 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_102,_zz_sbuf_wdat_12_103}}}};
  assign _zz_sbuf_wdat_12_8 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_9 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_10,_zz_sbuf_wdat_12_11}}}};
  assign _zz_sbuf_wdat_12_40 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_41 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_42,_zz_sbuf_wdat_12_43}}}};
  assign _zz_sbuf_wdat_12_72 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_73 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_74,_zz_sbuf_wdat_12_75}}}};
  assign _zz_sbuf_wdat_12_102 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_103 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_104,_zz_sbuf_wdat_12_105}}}};
  assign _zz_sbuf_wdat_12_10 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_11 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_12,_zz_sbuf_wdat_12_13}}}};
  assign _zz_sbuf_wdat_12_42 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_43 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_44,_zz_sbuf_wdat_12_45}}}};
  assign _zz_sbuf_wdat_12_74 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_75 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_76,_zz_sbuf_wdat_12_77}}}};
  assign _zz_sbuf_wdat_12_104 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_105 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_106,_zz_sbuf_wdat_12_107}}}};
  assign _zz_sbuf_wdat_12_12 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_13 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_14,_zz_sbuf_wdat_12_15}}}};
  assign _zz_sbuf_wdat_12_44 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_45 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_46,_zz_sbuf_wdat_12_47}}}};
  assign _zz_sbuf_wdat_12_76 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_77 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_78,_zz_sbuf_wdat_12_79}}}};
  assign _zz_sbuf_wdat_12_106 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_107 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_108,_zz_sbuf_wdat_12_109}}}};
  assign _zz_sbuf_wdat_12_14 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_15 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_16,_zz_sbuf_wdat_12_17}}}};
  assign _zz_sbuf_wdat_12_46 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_47 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_48,_zz_sbuf_wdat_12_49}}}};
  assign _zz_sbuf_wdat_12_78 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_79 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_80,_zz_sbuf_wdat_12_81}}}};
  assign _zz_sbuf_wdat_12_108 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_109 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_110,_zz_sbuf_wdat_12_111}}}};
  assign _zz_sbuf_wdat_12_16 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_17 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_18,_zz_sbuf_wdat_12_19}}}};
  assign _zz_sbuf_wdat_12_48 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_49 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_50,_zz_sbuf_wdat_12_51}}}};
  assign _zz_sbuf_wdat_12_80 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_81 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_82,_zz_sbuf_wdat_12_83}}}};
  assign _zz_sbuf_wdat_12_110 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_111 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_112,_zz_sbuf_wdat_12_113}}}};
  assign _zz_sbuf_wdat_12_18 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_19 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_20,_zz_sbuf_wdat_12_21}}}};
  assign _zz_sbuf_wdat_12_50 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_51 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_52,_zz_sbuf_wdat_12_53}}}};
  assign _zz_sbuf_wdat_12_82 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_83 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_84,_zz_sbuf_wdat_12_85}}}};
  assign _zz_sbuf_wdat_12_112 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_113 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_114,_zz_sbuf_wdat_12_115}}}};
  assign _zz_sbuf_wdat_12_20 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_21 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_22,_zz_sbuf_wdat_12_23}}}};
  assign _zz_sbuf_wdat_12_52 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_53 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_54,_zz_sbuf_wdat_12_55}}}};
  assign _zz_sbuf_wdat_12_84 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_85 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_86,_zz_sbuf_wdat_12_87}}}};
  assign _zz_sbuf_wdat_12_114 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_115 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_116,_zz_sbuf_wdat_12_117}}}};
  assign _zz_sbuf_wdat_12_22 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_23 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_24,_zz_sbuf_wdat_12_25}}}};
  assign _zz_sbuf_wdat_12_54 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_55 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_56,_zz_sbuf_wdat_12_57}}}};
  assign _zz_sbuf_wdat_12_86 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_87 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_88,_zz_sbuf_wdat_12_89}}}};
  assign _zz_sbuf_wdat_12_116 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_117 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_118,_zz_sbuf_wdat_12_119}}}};
  assign _zz_sbuf_wdat_12_24 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_25 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_26,_zz_sbuf_wdat_12_27}}}};
  assign _zz_sbuf_wdat_12_56 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_57 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_58,_zz_sbuf_wdat_12_59}}}};
  assign _zz_sbuf_wdat_12_88 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_89 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_90,_zz_sbuf_wdat_12_91}}}};
  assign _zz_sbuf_wdat_12_118 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_119 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_120,_zz_sbuf_wdat_12_121}}}};
  assign _zz_sbuf_wdat_12_26 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_27 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_28,_zz_sbuf_wdat_12_29}}}};
  assign _zz_sbuf_wdat_12_58 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_59 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_60,_zz_sbuf_wdat_12_61}}}};
  assign _zz_sbuf_wdat_12_90 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_91 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_92,_zz_sbuf_wdat_12_93}}}};
  assign _zz_sbuf_wdat_12_120 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_121 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_122,_zz_sbuf_wdat_12_123}}}};
  assign _zz_sbuf_wdat_12_28 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_29 = {dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_30,_zz_sbuf_wdat_12_31}}}}};
  assign _zz_sbuf_wdat_12_60 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_61 = {dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_62,_zz_sbuf_wdat_12_63}}}}};
  assign _zz_sbuf_wdat_12_92 = img2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_93 = {img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,img2sbuf_p0_wr_sel_12}}}};
  assign _zz_sbuf_wdat_12_122 = img2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_123 = {img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,img2sbuf_p1_wr_sel_12}}};
  assign _zz_sbuf_wdat_12_30 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_31 = dc2sbuf_p0_wr_sel_12;
  assign _zz_sbuf_wdat_12_62 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_12_63 = dc2sbuf_p1_wr_sel_12;
  assign _zz_sbuf_wdat_13 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_1 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_2,_zz_sbuf_wdat_13_3}}}};
  assign _zz_sbuf_wdat_13_32 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_33 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_34,_zz_sbuf_wdat_13_35}}}};
  assign _zz_sbuf_wdat_13_64 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_65 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_66,_zz_sbuf_wdat_13_67}}}};
  assign _zz_sbuf_wdat_13_94 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_95 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_96,_zz_sbuf_wdat_13_97}}}};
  assign _zz_sbuf_wdat_13_2 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_3 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_4,_zz_sbuf_wdat_13_5}}}};
  assign _zz_sbuf_wdat_13_34 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_35 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_36,_zz_sbuf_wdat_13_37}}}};
  assign _zz_sbuf_wdat_13_66 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_67 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_68,_zz_sbuf_wdat_13_69}}}};
  assign _zz_sbuf_wdat_13_96 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_97 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_98,_zz_sbuf_wdat_13_99}}}};
  assign _zz_sbuf_wdat_13_4 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_5 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_6,_zz_sbuf_wdat_13_7}}}};
  assign _zz_sbuf_wdat_13_36 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_37 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_38,_zz_sbuf_wdat_13_39}}}};
  assign _zz_sbuf_wdat_13_68 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_69 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_70,_zz_sbuf_wdat_13_71}}}};
  assign _zz_sbuf_wdat_13_98 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_99 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_100,_zz_sbuf_wdat_13_101}}}};
  assign _zz_sbuf_wdat_13_6 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_7 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_8,_zz_sbuf_wdat_13_9}}}};
  assign _zz_sbuf_wdat_13_38 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_39 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_40,_zz_sbuf_wdat_13_41}}}};
  assign _zz_sbuf_wdat_13_70 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_71 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_72,_zz_sbuf_wdat_13_73}}}};
  assign _zz_sbuf_wdat_13_100 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_101 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_102,_zz_sbuf_wdat_13_103}}}};
  assign _zz_sbuf_wdat_13_8 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_9 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_10,_zz_sbuf_wdat_13_11}}}};
  assign _zz_sbuf_wdat_13_40 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_41 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_42,_zz_sbuf_wdat_13_43}}}};
  assign _zz_sbuf_wdat_13_72 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_73 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_74,_zz_sbuf_wdat_13_75}}}};
  assign _zz_sbuf_wdat_13_102 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_103 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_104,_zz_sbuf_wdat_13_105}}}};
  assign _zz_sbuf_wdat_13_10 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_11 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_12,_zz_sbuf_wdat_13_13}}}};
  assign _zz_sbuf_wdat_13_42 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_43 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_44,_zz_sbuf_wdat_13_45}}}};
  assign _zz_sbuf_wdat_13_74 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_75 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_76,_zz_sbuf_wdat_13_77}}}};
  assign _zz_sbuf_wdat_13_104 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_105 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_106,_zz_sbuf_wdat_13_107}}}};
  assign _zz_sbuf_wdat_13_12 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_13 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_14,_zz_sbuf_wdat_13_15}}}};
  assign _zz_sbuf_wdat_13_44 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_45 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_46,_zz_sbuf_wdat_13_47}}}};
  assign _zz_sbuf_wdat_13_76 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_77 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_78,_zz_sbuf_wdat_13_79}}}};
  assign _zz_sbuf_wdat_13_106 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_107 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_108,_zz_sbuf_wdat_13_109}}}};
  assign _zz_sbuf_wdat_13_14 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_15 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_16,_zz_sbuf_wdat_13_17}}}};
  assign _zz_sbuf_wdat_13_46 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_47 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_48,_zz_sbuf_wdat_13_49}}}};
  assign _zz_sbuf_wdat_13_78 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_79 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_80,_zz_sbuf_wdat_13_81}}}};
  assign _zz_sbuf_wdat_13_108 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_109 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_110,_zz_sbuf_wdat_13_111}}}};
  assign _zz_sbuf_wdat_13_16 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_17 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_18,_zz_sbuf_wdat_13_19}}}};
  assign _zz_sbuf_wdat_13_48 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_49 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_50,_zz_sbuf_wdat_13_51}}}};
  assign _zz_sbuf_wdat_13_80 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_81 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_82,_zz_sbuf_wdat_13_83}}}};
  assign _zz_sbuf_wdat_13_110 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_111 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_112,_zz_sbuf_wdat_13_113}}}};
  assign _zz_sbuf_wdat_13_18 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_19 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_20,_zz_sbuf_wdat_13_21}}}};
  assign _zz_sbuf_wdat_13_50 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_51 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_52,_zz_sbuf_wdat_13_53}}}};
  assign _zz_sbuf_wdat_13_82 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_83 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_84,_zz_sbuf_wdat_13_85}}}};
  assign _zz_sbuf_wdat_13_112 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_113 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_114,_zz_sbuf_wdat_13_115}}}};
  assign _zz_sbuf_wdat_13_20 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_21 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_22,_zz_sbuf_wdat_13_23}}}};
  assign _zz_sbuf_wdat_13_52 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_53 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_54,_zz_sbuf_wdat_13_55}}}};
  assign _zz_sbuf_wdat_13_84 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_85 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_86,_zz_sbuf_wdat_13_87}}}};
  assign _zz_sbuf_wdat_13_114 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_115 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_116,_zz_sbuf_wdat_13_117}}}};
  assign _zz_sbuf_wdat_13_22 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_23 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_24,_zz_sbuf_wdat_13_25}}}};
  assign _zz_sbuf_wdat_13_54 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_55 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_56,_zz_sbuf_wdat_13_57}}}};
  assign _zz_sbuf_wdat_13_86 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_87 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_88,_zz_sbuf_wdat_13_89}}}};
  assign _zz_sbuf_wdat_13_116 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_117 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_118,_zz_sbuf_wdat_13_119}}}};
  assign _zz_sbuf_wdat_13_24 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_25 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_26,_zz_sbuf_wdat_13_27}}}};
  assign _zz_sbuf_wdat_13_56 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_57 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_58,_zz_sbuf_wdat_13_59}}}};
  assign _zz_sbuf_wdat_13_88 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_89 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_90,_zz_sbuf_wdat_13_91}}}};
  assign _zz_sbuf_wdat_13_118 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_119 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_120,_zz_sbuf_wdat_13_121}}}};
  assign _zz_sbuf_wdat_13_26 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_27 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_28,_zz_sbuf_wdat_13_29}}}};
  assign _zz_sbuf_wdat_13_58 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_59 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_60,_zz_sbuf_wdat_13_61}}}};
  assign _zz_sbuf_wdat_13_90 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_91 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_92,_zz_sbuf_wdat_13_93}}}};
  assign _zz_sbuf_wdat_13_120 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_121 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_122,_zz_sbuf_wdat_13_123}}}};
  assign _zz_sbuf_wdat_13_28 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_29 = {dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_30,_zz_sbuf_wdat_13_31}}}}};
  assign _zz_sbuf_wdat_13_60 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_61 = {dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_62,_zz_sbuf_wdat_13_63}}}}};
  assign _zz_sbuf_wdat_13_92 = img2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_93 = {img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,img2sbuf_p0_wr_sel_13}}}};
  assign _zz_sbuf_wdat_13_122 = img2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_123 = {img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,img2sbuf_p1_wr_sel_13}}};
  assign _zz_sbuf_wdat_13_30 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_31 = dc2sbuf_p0_wr_sel_13;
  assign _zz_sbuf_wdat_13_62 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_13_63 = dc2sbuf_p1_wr_sel_13;
  assign _zz_sbuf_wdat_14 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_1 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_2,_zz_sbuf_wdat_14_3}}}};
  assign _zz_sbuf_wdat_14_32 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_33 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_34,_zz_sbuf_wdat_14_35}}}};
  assign _zz_sbuf_wdat_14_64 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_65 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_66,_zz_sbuf_wdat_14_67}}}};
  assign _zz_sbuf_wdat_14_94 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_95 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_96,_zz_sbuf_wdat_14_97}}}};
  assign _zz_sbuf_wdat_14_2 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_3 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_4,_zz_sbuf_wdat_14_5}}}};
  assign _zz_sbuf_wdat_14_34 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_35 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_36,_zz_sbuf_wdat_14_37}}}};
  assign _zz_sbuf_wdat_14_66 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_67 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_68,_zz_sbuf_wdat_14_69}}}};
  assign _zz_sbuf_wdat_14_96 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_97 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_98,_zz_sbuf_wdat_14_99}}}};
  assign _zz_sbuf_wdat_14_4 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_5 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_6,_zz_sbuf_wdat_14_7}}}};
  assign _zz_sbuf_wdat_14_36 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_37 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_38,_zz_sbuf_wdat_14_39}}}};
  assign _zz_sbuf_wdat_14_68 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_69 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_70,_zz_sbuf_wdat_14_71}}}};
  assign _zz_sbuf_wdat_14_98 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_99 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_100,_zz_sbuf_wdat_14_101}}}};
  assign _zz_sbuf_wdat_14_6 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_7 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_8,_zz_sbuf_wdat_14_9}}}};
  assign _zz_sbuf_wdat_14_38 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_39 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_40,_zz_sbuf_wdat_14_41}}}};
  assign _zz_sbuf_wdat_14_70 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_71 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_72,_zz_sbuf_wdat_14_73}}}};
  assign _zz_sbuf_wdat_14_100 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_101 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_102,_zz_sbuf_wdat_14_103}}}};
  assign _zz_sbuf_wdat_14_8 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_9 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_10,_zz_sbuf_wdat_14_11}}}};
  assign _zz_sbuf_wdat_14_40 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_41 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_42,_zz_sbuf_wdat_14_43}}}};
  assign _zz_sbuf_wdat_14_72 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_73 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_74,_zz_sbuf_wdat_14_75}}}};
  assign _zz_sbuf_wdat_14_102 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_103 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_104,_zz_sbuf_wdat_14_105}}}};
  assign _zz_sbuf_wdat_14_10 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_11 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_12,_zz_sbuf_wdat_14_13}}}};
  assign _zz_sbuf_wdat_14_42 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_43 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_44,_zz_sbuf_wdat_14_45}}}};
  assign _zz_sbuf_wdat_14_74 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_75 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_76,_zz_sbuf_wdat_14_77}}}};
  assign _zz_sbuf_wdat_14_104 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_105 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_106,_zz_sbuf_wdat_14_107}}}};
  assign _zz_sbuf_wdat_14_12 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_13 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_14,_zz_sbuf_wdat_14_15}}}};
  assign _zz_sbuf_wdat_14_44 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_45 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_46,_zz_sbuf_wdat_14_47}}}};
  assign _zz_sbuf_wdat_14_76 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_77 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_78,_zz_sbuf_wdat_14_79}}}};
  assign _zz_sbuf_wdat_14_106 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_107 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_108,_zz_sbuf_wdat_14_109}}}};
  assign _zz_sbuf_wdat_14_14 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_15 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_16,_zz_sbuf_wdat_14_17}}}};
  assign _zz_sbuf_wdat_14_46 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_47 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_48,_zz_sbuf_wdat_14_49}}}};
  assign _zz_sbuf_wdat_14_78 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_79 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_80,_zz_sbuf_wdat_14_81}}}};
  assign _zz_sbuf_wdat_14_108 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_109 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_110,_zz_sbuf_wdat_14_111}}}};
  assign _zz_sbuf_wdat_14_16 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_17 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_18,_zz_sbuf_wdat_14_19}}}};
  assign _zz_sbuf_wdat_14_48 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_49 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_50,_zz_sbuf_wdat_14_51}}}};
  assign _zz_sbuf_wdat_14_80 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_81 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_82,_zz_sbuf_wdat_14_83}}}};
  assign _zz_sbuf_wdat_14_110 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_111 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_112,_zz_sbuf_wdat_14_113}}}};
  assign _zz_sbuf_wdat_14_18 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_19 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_20,_zz_sbuf_wdat_14_21}}}};
  assign _zz_sbuf_wdat_14_50 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_51 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_52,_zz_sbuf_wdat_14_53}}}};
  assign _zz_sbuf_wdat_14_82 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_83 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_84,_zz_sbuf_wdat_14_85}}}};
  assign _zz_sbuf_wdat_14_112 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_113 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_114,_zz_sbuf_wdat_14_115}}}};
  assign _zz_sbuf_wdat_14_20 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_21 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_22,_zz_sbuf_wdat_14_23}}}};
  assign _zz_sbuf_wdat_14_52 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_53 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_54,_zz_sbuf_wdat_14_55}}}};
  assign _zz_sbuf_wdat_14_84 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_85 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_86,_zz_sbuf_wdat_14_87}}}};
  assign _zz_sbuf_wdat_14_114 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_115 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_116,_zz_sbuf_wdat_14_117}}}};
  assign _zz_sbuf_wdat_14_22 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_23 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_24,_zz_sbuf_wdat_14_25}}}};
  assign _zz_sbuf_wdat_14_54 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_55 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_56,_zz_sbuf_wdat_14_57}}}};
  assign _zz_sbuf_wdat_14_86 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_87 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_88,_zz_sbuf_wdat_14_89}}}};
  assign _zz_sbuf_wdat_14_116 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_117 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_118,_zz_sbuf_wdat_14_119}}}};
  assign _zz_sbuf_wdat_14_24 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_25 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_26,_zz_sbuf_wdat_14_27}}}};
  assign _zz_sbuf_wdat_14_56 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_57 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_58,_zz_sbuf_wdat_14_59}}}};
  assign _zz_sbuf_wdat_14_88 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_89 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_90,_zz_sbuf_wdat_14_91}}}};
  assign _zz_sbuf_wdat_14_118 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_119 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_120,_zz_sbuf_wdat_14_121}}}};
  assign _zz_sbuf_wdat_14_26 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_27 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_28,_zz_sbuf_wdat_14_29}}}};
  assign _zz_sbuf_wdat_14_58 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_59 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_60,_zz_sbuf_wdat_14_61}}}};
  assign _zz_sbuf_wdat_14_90 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_91 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_92,_zz_sbuf_wdat_14_93}}}};
  assign _zz_sbuf_wdat_14_120 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_121 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_122,_zz_sbuf_wdat_14_123}}}};
  assign _zz_sbuf_wdat_14_28 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_29 = {dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_30,_zz_sbuf_wdat_14_31}}}}};
  assign _zz_sbuf_wdat_14_60 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_61 = {dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_62,_zz_sbuf_wdat_14_63}}}}};
  assign _zz_sbuf_wdat_14_92 = img2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_93 = {img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,img2sbuf_p0_wr_sel_14}}}};
  assign _zz_sbuf_wdat_14_122 = img2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_123 = {img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,img2sbuf_p1_wr_sel_14}}};
  assign _zz_sbuf_wdat_14_30 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_31 = dc2sbuf_p0_wr_sel_14;
  assign _zz_sbuf_wdat_14_62 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_14_63 = dc2sbuf_p1_wr_sel_14;
  assign _zz_sbuf_wdat_15 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_1 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_2,_zz_sbuf_wdat_15_3}}}};
  assign _zz_sbuf_wdat_15_32 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_33 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_34,_zz_sbuf_wdat_15_35}}}};
  assign _zz_sbuf_wdat_15_64 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_65 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_66,_zz_sbuf_wdat_15_67}}}};
  assign _zz_sbuf_wdat_15_94 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_95 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_96,_zz_sbuf_wdat_15_97}}}};
  assign _zz_sbuf_wdat_15_2 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_3 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_4,_zz_sbuf_wdat_15_5}}}};
  assign _zz_sbuf_wdat_15_34 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_35 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_36,_zz_sbuf_wdat_15_37}}}};
  assign _zz_sbuf_wdat_15_66 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_67 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_68,_zz_sbuf_wdat_15_69}}}};
  assign _zz_sbuf_wdat_15_96 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_97 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_98,_zz_sbuf_wdat_15_99}}}};
  assign _zz_sbuf_wdat_15_4 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_5 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_6,_zz_sbuf_wdat_15_7}}}};
  assign _zz_sbuf_wdat_15_36 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_37 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_38,_zz_sbuf_wdat_15_39}}}};
  assign _zz_sbuf_wdat_15_68 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_69 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_70,_zz_sbuf_wdat_15_71}}}};
  assign _zz_sbuf_wdat_15_98 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_99 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_100,_zz_sbuf_wdat_15_101}}}};
  assign _zz_sbuf_wdat_15_6 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_7 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_8,_zz_sbuf_wdat_15_9}}}};
  assign _zz_sbuf_wdat_15_38 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_39 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_40,_zz_sbuf_wdat_15_41}}}};
  assign _zz_sbuf_wdat_15_70 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_71 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_72,_zz_sbuf_wdat_15_73}}}};
  assign _zz_sbuf_wdat_15_100 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_101 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_102,_zz_sbuf_wdat_15_103}}}};
  assign _zz_sbuf_wdat_15_8 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_9 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_10,_zz_sbuf_wdat_15_11}}}};
  assign _zz_sbuf_wdat_15_40 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_41 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_42,_zz_sbuf_wdat_15_43}}}};
  assign _zz_sbuf_wdat_15_72 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_73 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_74,_zz_sbuf_wdat_15_75}}}};
  assign _zz_sbuf_wdat_15_102 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_103 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_104,_zz_sbuf_wdat_15_105}}}};
  assign _zz_sbuf_wdat_15_10 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_11 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_12,_zz_sbuf_wdat_15_13}}}};
  assign _zz_sbuf_wdat_15_42 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_43 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_44,_zz_sbuf_wdat_15_45}}}};
  assign _zz_sbuf_wdat_15_74 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_75 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_76,_zz_sbuf_wdat_15_77}}}};
  assign _zz_sbuf_wdat_15_104 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_105 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_106,_zz_sbuf_wdat_15_107}}}};
  assign _zz_sbuf_wdat_15_12 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_13 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_14,_zz_sbuf_wdat_15_15}}}};
  assign _zz_sbuf_wdat_15_44 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_45 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_46,_zz_sbuf_wdat_15_47}}}};
  assign _zz_sbuf_wdat_15_76 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_77 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_78,_zz_sbuf_wdat_15_79}}}};
  assign _zz_sbuf_wdat_15_106 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_107 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_108,_zz_sbuf_wdat_15_109}}}};
  assign _zz_sbuf_wdat_15_14 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_15 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_16,_zz_sbuf_wdat_15_17}}}};
  assign _zz_sbuf_wdat_15_46 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_47 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_48,_zz_sbuf_wdat_15_49}}}};
  assign _zz_sbuf_wdat_15_78 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_79 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_80,_zz_sbuf_wdat_15_81}}}};
  assign _zz_sbuf_wdat_15_108 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_109 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_110,_zz_sbuf_wdat_15_111}}}};
  assign _zz_sbuf_wdat_15_16 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_17 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_18,_zz_sbuf_wdat_15_19}}}};
  assign _zz_sbuf_wdat_15_48 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_49 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_50,_zz_sbuf_wdat_15_51}}}};
  assign _zz_sbuf_wdat_15_80 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_81 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_82,_zz_sbuf_wdat_15_83}}}};
  assign _zz_sbuf_wdat_15_110 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_111 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_112,_zz_sbuf_wdat_15_113}}}};
  assign _zz_sbuf_wdat_15_18 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_19 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_20,_zz_sbuf_wdat_15_21}}}};
  assign _zz_sbuf_wdat_15_50 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_51 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_52,_zz_sbuf_wdat_15_53}}}};
  assign _zz_sbuf_wdat_15_82 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_83 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_84,_zz_sbuf_wdat_15_85}}}};
  assign _zz_sbuf_wdat_15_112 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_113 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_114,_zz_sbuf_wdat_15_115}}}};
  assign _zz_sbuf_wdat_15_20 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_21 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_22,_zz_sbuf_wdat_15_23}}}};
  assign _zz_sbuf_wdat_15_52 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_53 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_54,_zz_sbuf_wdat_15_55}}}};
  assign _zz_sbuf_wdat_15_84 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_85 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_86,_zz_sbuf_wdat_15_87}}}};
  assign _zz_sbuf_wdat_15_114 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_115 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_116,_zz_sbuf_wdat_15_117}}}};
  assign _zz_sbuf_wdat_15_22 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_23 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_24,_zz_sbuf_wdat_15_25}}}};
  assign _zz_sbuf_wdat_15_54 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_55 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_56,_zz_sbuf_wdat_15_57}}}};
  assign _zz_sbuf_wdat_15_86 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_87 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_88,_zz_sbuf_wdat_15_89}}}};
  assign _zz_sbuf_wdat_15_116 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_117 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_118,_zz_sbuf_wdat_15_119}}}};
  assign _zz_sbuf_wdat_15_24 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_25 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_26,_zz_sbuf_wdat_15_27}}}};
  assign _zz_sbuf_wdat_15_56 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_57 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_58,_zz_sbuf_wdat_15_59}}}};
  assign _zz_sbuf_wdat_15_88 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_89 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_90,_zz_sbuf_wdat_15_91}}}};
  assign _zz_sbuf_wdat_15_118 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_119 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_120,_zz_sbuf_wdat_15_121}}}};
  assign _zz_sbuf_wdat_15_26 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_27 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_28,_zz_sbuf_wdat_15_29}}}};
  assign _zz_sbuf_wdat_15_58 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_59 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_60,_zz_sbuf_wdat_15_61}}}};
  assign _zz_sbuf_wdat_15_90 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_91 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_92,_zz_sbuf_wdat_15_93}}}};
  assign _zz_sbuf_wdat_15_120 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_121 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_122,_zz_sbuf_wdat_15_123}}}};
  assign _zz_sbuf_wdat_15_28 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_29 = {dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_30,_zz_sbuf_wdat_15_31}}}}};
  assign _zz_sbuf_wdat_15_60 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_61 = {dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_62,_zz_sbuf_wdat_15_63}}}}};
  assign _zz_sbuf_wdat_15_92 = img2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_93 = {img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,img2sbuf_p0_wr_sel_15}}}};
  assign _zz_sbuf_wdat_15_122 = img2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_123 = {img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,img2sbuf_p1_wr_sel_15}}};
  assign _zz_sbuf_wdat_15_30 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_31 = dc2sbuf_p0_wr_sel_15;
  assign _zz_sbuf_wdat_15_62 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_wdat_15_63 = dc2sbuf_p1_wr_sel_15;
  assign _zz_sbuf_ra_0 = dc2sbuf_p0_rd_sel_0;
  assign _zz_sbuf_ra_0_1 = {dc2sbuf_p0_rd_sel_0,{dc2sbuf_p0_rd_sel_0,dc2sbuf_p0_rd_sel_0}};
  assign _zz_sbuf_ra_0_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_0_3 = dc2sbuf_p1_rd_sel_0;
  assign _zz_sbuf_ra_0_4 = {dc2sbuf_p1_rd_sel_0,{dc2sbuf_p1_rd_sel_0,dc2sbuf_p1_rd_sel_0}};
  assign _zz_sbuf_ra_0_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_0_6 = img2sbuf_p0_rd_sel_0;
  assign _zz_sbuf_ra_0_7 = {img2sbuf_p0_rd_sel_0,img2sbuf_p0_rd_sel_0};
  assign _zz_sbuf_ra_0_8 = img2sbuf_p1_rd_sel_0;
  assign _zz_sbuf_ra_0_9 = img2sbuf_p1_rd_sel_0;
  assign _zz_sbuf_ra_1 = dc2sbuf_p0_rd_sel_1;
  assign _zz_sbuf_ra_1_1 = {dc2sbuf_p0_rd_sel_1,{dc2sbuf_p0_rd_sel_1,dc2sbuf_p0_rd_sel_1}};
  assign _zz_sbuf_ra_1_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_1_3 = dc2sbuf_p1_rd_sel_1;
  assign _zz_sbuf_ra_1_4 = {dc2sbuf_p1_rd_sel_1,{dc2sbuf_p1_rd_sel_1,dc2sbuf_p1_rd_sel_1}};
  assign _zz_sbuf_ra_1_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_1_6 = img2sbuf_p0_rd_sel_1;
  assign _zz_sbuf_ra_1_7 = {img2sbuf_p0_rd_sel_1,img2sbuf_p0_rd_sel_1};
  assign _zz_sbuf_ra_1_8 = img2sbuf_p1_rd_sel_1;
  assign _zz_sbuf_ra_1_9 = img2sbuf_p1_rd_sel_1;
  assign _zz_sbuf_ra_2 = dc2sbuf_p0_rd_sel_2;
  assign _zz_sbuf_ra_2_1 = {dc2sbuf_p0_rd_sel_2,{dc2sbuf_p0_rd_sel_2,dc2sbuf_p0_rd_sel_2}};
  assign _zz_sbuf_ra_2_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_2_3 = dc2sbuf_p1_rd_sel_2;
  assign _zz_sbuf_ra_2_4 = {dc2sbuf_p1_rd_sel_2,{dc2sbuf_p1_rd_sel_2,dc2sbuf_p1_rd_sel_2}};
  assign _zz_sbuf_ra_2_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_2_6 = img2sbuf_p0_rd_sel_2;
  assign _zz_sbuf_ra_2_7 = {img2sbuf_p0_rd_sel_2,img2sbuf_p0_rd_sel_2};
  assign _zz_sbuf_ra_2_8 = img2sbuf_p1_rd_sel_2;
  assign _zz_sbuf_ra_2_9 = img2sbuf_p1_rd_sel_2;
  assign _zz_sbuf_ra_3 = dc2sbuf_p0_rd_sel_3;
  assign _zz_sbuf_ra_3_1 = {dc2sbuf_p0_rd_sel_3,{dc2sbuf_p0_rd_sel_3,dc2sbuf_p0_rd_sel_3}};
  assign _zz_sbuf_ra_3_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_3_3 = dc2sbuf_p1_rd_sel_3;
  assign _zz_sbuf_ra_3_4 = {dc2sbuf_p1_rd_sel_3,{dc2sbuf_p1_rd_sel_3,dc2sbuf_p1_rd_sel_3}};
  assign _zz_sbuf_ra_3_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_3_6 = img2sbuf_p0_rd_sel_3;
  assign _zz_sbuf_ra_3_7 = {img2sbuf_p0_rd_sel_3,img2sbuf_p0_rd_sel_3};
  assign _zz_sbuf_ra_3_8 = img2sbuf_p1_rd_sel_3;
  assign _zz_sbuf_ra_3_9 = img2sbuf_p1_rd_sel_3;
  assign _zz_sbuf_ra_4 = dc2sbuf_p0_rd_sel_4;
  assign _zz_sbuf_ra_4_1 = {dc2sbuf_p0_rd_sel_4,{dc2sbuf_p0_rd_sel_4,dc2sbuf_p0_rd_sel_4}};
  assign _zz_sbuf_ra_4_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_4_3 = dc2sbuf_p1_rd_sel_4;
  assign _zz_sbuf_ra_4_4 = {dc2sbuf_p1_rd_sel_4,{dc2sbuf_p1_rd_sel_4,dc2sbuf_p1_rd_sel_4}};
  assign _zz_sbuf_ra_4_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_4_6 = img2sbuf_p0_rd_sel_4;
  assign _zz_sbuf_ra_4_7 = {img2sbuf_p0_rd_sel_4,img2sbuf_p0_rd_sel_4};
  assign _zz_sbuf_ra_4_8 = img2sbuf_p1_rd_sel_4;
  assign _zz_sbuf_ra_4_9 = img2sbuf_p1_rd_sel_4;
  assign _zz_sbuf_ra_5 = dc2sbuf_p0_rd_sel_5;
  assign _zz_sbuf_ra_5_1 = {dc2sbuf_p0_rd_sel_5,{dc2sbuf_p0_rd_sel_5,dc2sbuf_p0_rd_sel_5}};
  assign _zz_sbuf_ra_5_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_5_3 = dc2sbuf_p1_rd_sel_5;
  assign _zz_sbuf_ra_5_4 = {dc2sbuf_p1_rd_sel_5,{dc2sbuf_p1_rd_sel_5,dc2sbuf_p1_rd_sel_5}};
  assign _zz_sbuf_ra_5_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_5_6 = img2sbuf_p0_rd_sel_5;
  assign _zz_sbuf_ra_5_7 = {img2sbuf_p0_rd_sel_5,img2sbuf_p0_rd_sel_5};
  assign _zz_sbuf_ra_5_8 = img2sbuf_p1_rd_sel_5;
  assign _zz_sbuf_ra_5_9 = img2sbuf_p1_rd_sel_5;
  assign _zz_sbuf_ra_6 = dc2sbuf_p0_rd_sel_6;
  assign _zz_sbuf_ra_6_1 = {dc2sbuf_p0_rd_sel_6,{dc2sbuf_p0_rd_sel_6,dc2sbuf_p0_rd_sel_6}};
  assign _zz_sbuf_ra_6_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_6_3 = dc2sbuf_p1_rd_sel_6;
  assign _zz_sbuf_ra_6_4 = {dc2sbuf_p1_rd_sel_6,{dc2sbuf_p1_rd_sel_6,dc2sbuf_p1_rd_sel_6}};
  assign _zz_sbuf_ra_6_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_6_6 = img2sbuf_p0_rd_sel_6;
  assign _zz_sbuf_ra_6_7 = {img2sbuf_p0_rd_sel_6,img2sbuf_p0_rd_sel_6};
  assign _zz_sbuf_ra_6_8 = img2sbuf_p1_rd_sel_6;
  assign _zz_sbuf_ra_6_9 = img2sbuf_p1_rd_sel_6;
  assign _zz_sbuf_ra_7 = dc2sbuf_p0_rd_sel_7;
  assign _zz_sbuf_ra_7_1 = {dc2sbuf_p0_rd_sel_7,{dc2sbuf_p0_rd_sel_7,dc2sbuf_p0_rd_sel_7}};
  assign _zz_sbuf_ra_7_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_7_3 = dc2sbuf_p1_rd_sel_7;
  assign _zz_sbuf_ra_7_4 = {dc2sbuf_p1_rd_sel_7,{dc2sbuf_p1_rd_sel_7,dc2sbuf_p1_rd_sel_7}};
  assign _zz_sbuf_ra_7_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_7_6 = img2sbuf_p0_rd_sel_7;
  assign _zz_sbuf_ra_7_7 = {img2sbuf_p0_rd_sel_7,img2sbuf_p0_rd_sel_7};
  assign _zz_sbuf_ra_7_8 = img2sbuf_p1_rd_sel_7;
  assign _zz_sbuf_ra_7_9 = img2sbuf_p1_rd_sel_7;
  assign _zz_sbuf_ra_8 = dc2sbuf_p0_rd_sel_8;
  assign _zz_sbuf_ra_8_1 = {dc2sbuf_p0_rd_sel_8,{dc2sbuf_p0_rd_sel_8,dc2sbuf_p0_rd_sel_8}};
  assign _zz_sbuf_ra_8_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_8_3 = dc2sbuf_p1_rd_sel_8;
  assign _zz_sbuf_ra_8_4 = {dc2sbuf_p1_rd_sel_8,{dc2sbuf_p1_rd_sel_8,dc2sbuf_p1_rd_sel_8}};
  assign _zz_sbuf_ra_8_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_8_6 = img2sbuf_p0_rd_sel_8;
  assign _zz_sbuf_ra_8_7 = {img2sbuf_p0_rd_sel_8,img2sbuf_p0_rd_sel_8};
  assign _zz_sbuf_ra_8_8 = img2sbuf_p1_rd_sel_8;
  assign _zz_sbuf_ra_8_9 = img2sbuf_p1_rd_sel_8;
  assign _zz_sbuf_ra_9 = dc2sbuf_p0_rd_sel_9;
  assign _zz_sbuf_ra_9_1 = {dc2sbuf_p0_rd_sel_9,{dc2sbuf_p0_rd_sel_9,dc2sbuf_p0_rd_sel_9}};
  assign _zz_sbuf_ra_9_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_9_3 = dc2sbuf_p1_rd_sel_9;
  assign _zz_sbuf_ra_9_4 = {dc2sbuf_p1_rd_sel_9,{dc2sbuf_p1_rd_sel_9,dc2sbuf_p1_rd_sel_9}};
  assign _zz_sbuf_ra_9_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_9_6 = img2sbuf_p0_rd_sel_9;
  assign _zz_sbuf_ra_9_7 = {img2sbuf_p0_rd_sel_9,img2sbuf_p0_rd_sel_9};
  assign _zz_sbuf_ra_9_8 = img2sbuf_p1_rd_sel_9;
  assign _zz_sbuf_ra_9_9 = img2sbuf_p1_rd_sel_9;
  assign _zz_sbuf_ra_10 = dc2sbuf_p0_rd_sel_10;
  assign _zz_sbuf_ra_10_1 = {dc2sbuf_p0_rd_sel_10,{dc2sbuf_p0_rd_sel_10,dc2sbuf_p0_rd_sel_10}};
  assign _zz_sbuf_ra_10_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_10_3 = dc2sbuf_p1_rd_sel_10;
  assign _zz_sbuf_ra_10_4 = {dc2sbuf_p1_rd_sel_10,{dc2sbuf_p1_rd_sel_10,dc2sbuf_p1_rd_sel_10}};
  assign _zz_sbuf_ra_10_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_10_6 = img2sbuf_p0_rd_sel_10;
  assign _zz_sbuf_ra_10_7 = {img2sbuf_p0_rd_sel_10,img2sbuf_p0_rd_sel_10};
  assign _zz_sbuf_ra_10_8 = img2sbuf_p1_rd_sel_10;
  assign _zz_sbuf_ra_10_9 = img2sbuf_p1_rd_sel_10;
  assign _zz_sbuf_ra_11 = dc2sbuf_p0_rd_sel_11;
  assign _zz_sbuf_ra_11_1 = {dc2sbuf_p0_rd_sel_11,{dc2sbuf_p0_rd_sel_11,dc2sbuf_p0_rd_sel_11}};
  assign _zz_sbuf_ra_11_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_11_3 = dc2sbuf_p1_rd_sel_11;
  assign _zz_sbuf_ra_11_4 = {dc2sbuf_p1_rd_sel_11,{dc2sbuf_p1_rd_sel_11,dc2sbuf_p1_rd_sel_11}};
  assign _zz_sbuf_ra_11_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_11_6 = img2sbuf_p0_rd_sel_11;
  assign _zz_sbuf_ra_11_7 = {img2sbuf_p0_rd_sel_11,img2sbuf_p0_rd_sel_11};
  assign _zz_sbuf_ra_11_8 = img2sbuf_p1_rd_sel_11;
  assign _zz_sbuf_ra_11_9 = img2sbuf_p1_rd_sel_11;
  assign _zz_sbuf_ra_12 = dc2sbuf_p0_rd_sel_12;
  assign _zz_sbuf_ra_12_1 = {dc2sbuf_p0_rd_sel_12,{dc2sbuf_p0_rd_sel_12,dc2sbuf_p0_rd_sel_12}};
  assign _zz_sbuf_ra_12_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_12_3 = dc2sbuf_p1_rd_sel_12;
  assign _zz_sbuf_ra_12_4 = {dc2sbuf_p1_rd_sel_12,{dc2sbuf_p1_rd_sel_12,dc2sbuf_p1_rd_sel_12}};
  assign _zz_sbuf_ra_12_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_12_6 = img2sbuf_p0_rd_sel_12;
  assign _zz_sbuf_ra_12_7 = {img2sbuf_p0_rd_sel_12,img2sbuf_p0_rd_sel_12};
  assign _zz_sbuf_ra_12_8 = img2sbuf_p1_rd_sel_12;
  assign _zz_sbuf_ra_12_9 = img2sbuf_p1_rd_sel_12;
  assign _zz_sbuf_ra_13 = dc2sbuf_p0_rd_sel_13;
  assign _zz_sbuf_ra_13_1 = {dc2sbuf_p0_rd_sel_13,{dc2sbuf_p0_rd_sel_13,dc2sbuf_p0_rd_sel_13}};
  assign _zz_sbuf_ra_13_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_13_3 = dc2sbuf_p1_rd_sel_13;
  assign _zz_sbuf_ra_13_4 = {dc2sbuf_p1_rd_sel_13,{dc2sbuf_p1_rd_sel_13,dc2sbuf_p1_rd_sel_13}};
  assign _zz_sbuf_ra_13_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_13_6 = img2sbuf_p0_rd_sel_13;
  assign _zz_sbuf_ra_13_7 = {img2sbuf_p0_rd_sel_13,img2sbuf_p0_rd_sel_13};
  assign _zz_sbuf_ra_13_8 = img2sbuf_p1_rd_sel_13;
  assign _zz_sbuf_ra_13_9 = img2sbuf_p1_rd_sel_13;
  assign _zz_sbuf_ra_14 = dc2sbuf_p0_rd_sel_14;
  assign _zz_sbuf_ra_14_1 = {dc2sbuf_p0_rd_sel_14,{dc2sbuf_p0_rd_sel_14,dc2sbuf_p0_rd_sel_14}};
  assign _zz_sbuf_ra_14_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_14_3 = dc2sbuf_p1_rd_sel_14;
  assign _zz_sbuf_ra_14_4 = {dc2sbuf_p1_rd_sel_14,{dc2sbuf_p1_rd_sel_14,dc2sbuf_p1_rd_sel_14}};
  assign _zz_sbuf_ra_14_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_14_6 = img2sbuf_p0_rd_sel_14;
  assign _zz_sbuf_ra_14_7 = {img2sbuf_p0_rd_sel_14,img2sbuf_p0_rd_sel_14};
  assign _zz_sbuf_ra_14_8 = img2sbuf_p1_rd_sel_14;
  assign _zz_sbuf_ra_14_9 = img2sbuf_p1_rd_sel_14;
  assign _zz_sbuf_ra_15 = dc2sbuf_p0_rd_sel_15;
  assign _zz_sbuf_ra_15_1 = {dc2sbuf_p0_rd_sel_15,{dc2sbuf_p0_rd_sel_15,dc2sbuf_p0_rd_sel_15}};
  assign _zz_sbuf_ra_15_2 = dc2sbuf_p_rd_0_addr_payload[3 : 0];
  assign _zz_sbuf_ra_15_3 = dc2sbuf_p1_rd_sel_15;
  assign _zz_sbuf_ra_15_4 = {dc2sbuf_p1_rd_sel_15,{dc2sbuf_p1_rd_sel_15,dc2sbuf_p1_rd_sel_15}};
  assign _zz_sbuf_ra_15_5 = dc2sbuf_p_rd_1_addr_payload[3 : 0];
  assign _zz_sbuf_ra_15_6 = img2sbuf_p0_rd_sel_15;
  assign _zz_sbuf_ra_15_7 = {img2sbuf_p0_rd_sel_15,img2sbuf_p0_rd_sel_15};
  assign _zz_sbuf_ra_15_8 = img2sbuf_p1_rd_sel_15;
  assign _zz_sbuf_ra_15_9 = img2sbuf_p1_rd_sel_15;
  assign _zz_shareBuffer_sbuf_p0_rdat = (((_zz_shareBuffer_sbuf_p0_rdat_1 | _zz_shareBuffer_sbuf_p0_rdat_895) | (_zz_shareBuffer_sbuf_p0_rdat_1008 & shareBuffer_sbuf_rdat_9)) | ({_zz_shareBuffer_sbuf_p0_rdat_1121,_zz_shareBuffer_sbuf_p0_rdat_1122} & shareBuffer_sbuf_rdat_10));
  assign _zz_shareBuffer_sbuf_p0_rdat_1233 = ({shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1234,_zz_shareBuffer_sbuf_p0_rdat_1235}} & shareBuffer_sbuf_rdat_11);
  assign _zz_shareBuffer_sbuf_p0_rdat_1346 = {shareBuffer_sbuf_p0_re_norm_d1_12,{shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1347,_zz_shareBuffer_sbuf_p0_rdat_1348}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1457 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1458 = {shareBuffer_sbuf_p0_re_norm_d1_13,{shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1459,_zz_shareBuffer_sbuf_p0_rdat_1460}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1569 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1570 = {shareBuffer_sbuf_p0_re_norm_d1_14,{shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1571,_zz_shareBuffer_sbuf_p0_rdat_1572}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1679 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1680 = {shareBuffer_sbuf_p0_re_norm_d1_15,{shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1681,_zz_shareBuffer_sbuf_p0_rdat_1682}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1 = ((_zz_shareBuffer_sbuf_p0_rdat_2 | _zz_shareBuffer_sbuf_p0_rdat_669) | (_zz_shareBuffer_sbuf_p0_rdat_782 & shareBuffer_sbuf_rdat_7));
  assign _zz_shareBuffer_sbuf_p0_rdat_895 = ({_zz_shareBuffer_sbuf_p0_rdat_896,_zz_shareBuffer_sbuf_p0_rdat_897} & shareBuffer_sbuf_rdat_8);
  assign _zz_shareBuffer_sbuf_p0_rdat_1008 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1009,_zz_shareBuffer_sbuf_p0_rdat_1010}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1121 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1122 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1123,_zz_shareBuffer_sbuf_p0_rdat_1124}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1234 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1235 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1236,_zz_shareBuffer_sbuf_p0_rdat_1237}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1347 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1348 = {shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1349,_zz_shareBuffer_sbuf_p0_rdat_1350}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1459 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1460 = {shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1461,_zz_shareBuffer_sbuf_p0_rdat_1462}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1571 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1572 = {shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1573,_zz_shareBuffer_sbuf_p0_rdat_1574}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1681 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1682 = {shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1683,_zz_shareBuffer_sbuf_p0_rdat_1684}};
  assign _zz_shareBuffer_sbuf_p0_rdat_2 = ((_zz_shareBuffer_sbuf_p0_rdat_3 | _zz_shareBuffer_sbuf_p0_rdat_445) | (_zz_shareBuffer_sbuf_p0_rdat_558 & shareBuffer_sbuf_rdat_5));
  assign _zz_shareBuffer_sbuf_p0_rdat_669 = ({_zz_shareBuffer_sbuf_p0_rdat_670,_zz_shareBuffer_sbuf_p0_rdat_671} & shareBuffer_sbuf_rdat_6);
  assign _zz_shareBuffer_sbuf_p0_rdat_782 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_783,_zz_shareBuffer_sbuf_p0_rdat_784}};
  assign _zz_shareBuffer_sbuf_p0_rdat_896 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_897 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_898,_zz_shareBuffer_sbuf_p0_rdat_899}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1009 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1010 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1011,_zz_shareBuffer_sbuf_p0_rdat_1012}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1123 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1124 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1125,_zz_shareBuffer_sbuf_p0_rdat_1126}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1236 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1237 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1238,_zz_shareBuffer_sbuf_p0_rdat_1239}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1349 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1350 = {shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1351,_zz_shareBuffer_sbuf_p0_rdat_1352}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1461 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1462 = {shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1463,_zz_shareBuffer_sbuf_p0_rdat_1464}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1573 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1574 = {shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1575,_zz_shareBuffer_sbuf_p0_rdat_1576}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1683 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1684 = {shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1685,_zz_shareBuffer_sbuf_p0_rdat_1686}};
  assign _zz_shareBuffer_sbuf_p0_rdat_3 = ((_zz_shareBuffer_sbuf_p0_rdat_4 | _zz_shareBuffer_sbuf_p0_rdat_223) | (_zz_shareBuffer_sbuf_p0_rdat_334 & shareBuffer_sbuf_rdat_3));
  assign _zz_shareBuffer_sbuf_p0_rdat_445 = ({_zz_shareBuffer_sbuf_p0_rdat_446,_zz_shareBuffer_sbuf_p0_rdat_447} & shareBuffer_sbuf_rdat_4);
  assign _zz_shareBuffer_sbuf_p0_rdat_558 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_559,_zz_shareBuffer_sbuf_p0_rdat_560}};
  assign _zz_shareBuffer_sbuf_p0_rdat_670 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_671 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_672,_zz_shareBuffer_sbuf_p0_rdat_673}};
  assign _zz_shareBuffer_sbuf_p0_rdat_783 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_784 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_785,_zz_shareBuffer_sbuf_p0_rdat_786}};
  assign _zz_shareBuffer_sbuf_p0_rdat_898 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_899 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_900,_zz_shareBuffer_sbuf_p0_rdat_901}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1011 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1012 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1013,_zz_shareBuffer_sbuf_p0_rdat_1014}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1125 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1126 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1127,_zz_shareBuffer_sbuf_p0_rdat_1128}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1238 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1239 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1240,_zz_shareBuffer_sbuf_p0_rdat_1241}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1351 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1352 = {shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1353,_zz_shareBuffer_sbuf_p0_rdat_1354}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1463 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1464 = {shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1465,_zz_shareBuffer_sbuf_p0_rdat_1466}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1575 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1576 = {shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1577,_zz_shareBuffer_sbuf_p0_rdat_1578}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1685 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1686 = {shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1687,_zz_shareBuffer_sbuf_p0_rdat_1688}};
  assign _zz_shareBuffer_sbuf_p0_rdat_4 = ((_zz_shareBuffer_sbuf_p0_rdat_5 & shareBuffer_sbuf_rdat_0) | (_zz_shareBuffer_sbuf_p0_rdat_114 & shareBuffer_sbuf_rdat_1));
  assign _zz_shareBuffer_sbuf_p0_rdat_223 = ({_zz_shareBuffer_sbuf_p0_rdat_224,_zz_shareBuffer_sbuf_p0_rdat_225} & shareBuffer_sbuf_rdat_2);
  assign _zz_shareBuffer_sbuf_p0_rdat_334 = {shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_335,_zz_shareBuffer_sbuf_p0_rdat_336}};
  assign _zz_shareBuffer_sbuf_p0_rdat_446 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_447 = {shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_448,_zz_shareBuffer_sbuf_p0_rdat_449}};
  assign _zz_shareBuffer_sbuf_p0_rdat_559 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_560 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_561,_zz_shareBuffer_sbuf_p0_rdat_562}};
  assign _zz_shareBuffer_sbuf_p0_rdat_672 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_673 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_674,_zz_shareBuffer_sbuf_p0_rdat_675}};
  assign _zz_shareBuffer_sbuf_p0_rdat_785 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_786 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_787,_zz_shareBuffer_sbuf_p0_rdat_788}};
  assign _zz_shareBuffer_sbuf_p0_rdat_900 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_901 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_902,_zz_shareBuffer_sbuf_p0_rdat_903}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1013 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1014 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1015,_zz_shareBuffer_sbuf_p0_rdat_1016}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1127 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1128 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1129,_zz_shareBuffer_sbuf_p0_rdat_1130}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1240 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1241 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1242,_zz_shareBuffer_sbuf_p0_rdat_1243}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1353 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1354 = {shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1355,_zz_shareBuffer_sbuf_p0_rdat_1356}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1465 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1466 = {shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1467,_zz_shareBuffer_sbuf_p0_rdat_1468}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1577 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1578 = {shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1579,_zz_shareBuffer_sbuf_p0_rdat_1580}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1687 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1688 = {shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1689,_zz_shareBuffer_sbuf_p0_rdat_1690}};
  assign _zz_shareBuffer_sbuf_p0_rdat_5 = {_zz_shareBuffer_sbuf_p0_rdat_6,_zz_shareBuffer_sbuf_p0_rdat_7};
  assign _zz_shareBuffer_sbuf_p0_rdat_114 = {_zz_shareBuffer_sbuf_p0_rdat_115,_zz_shareBuffer_sbuf_p0_rdat_116};
  assign _zz_shareBuffer_sbuf_p0_rdat_224 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_225 = {_zz_shareBuffer_sbuf_p0_rdat_226,_zz_shareBuffer_sbuf_p0_rdat_227};
  assign _zz_shareBuffer_sbuf_p0_rdat_335 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_336 = {_zz_shareBuffer_sbuf_p0_rdat_337,_zz_shareBuffer_sbuf_p0_rdat_338};
  assign _zz_shareBuffer_sbuf_p0_rdat_448 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_449 = {_zz_shareBuffer_sbuf_p0_rdat_450,_zz_shareBuffer_sbuf_p0_rdat_451};
  assign _zz_shareBuffer_sbuf_p0_rdat_561 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_562 = {_zz_shareBuffer_sbuf_p0_rdat_563,_zz_shareBuffer_sbuf_p0_rdat_564};
  assign _zz_shareBuffer_sbuf_p0_rdat_674 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_675 = {_zz_shareBuffer_sbuf_p0_rdat_676,_zz_shareBuffer_sbuf_p0_rdat_677};
  assign _zz_shareBuffer_sbuf_p0_rdat_787 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_788 = {_zz_shareBuffer_sbuf_p0_rdat_789,_zz_shareBuffer_sbuf_p0_rdat_790};
  assign _zz_shareBuffer_sbuf_p0_rdat_902 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_903 = {_zz_shareBuffer_sbuf_p0_rdat_904,_zz_shareBuffer_sbuf_p0_rdat_905};
  assign _zz_shareBuffer_sbuf_p0_rdat_1015 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1016 = {_zz_shareBuffer_sbuf_p0_rdat_1017,_zz_shareBuffer_sbuf_p0_rdat_1018};
  assign _zz_shareBuffer_sbuf_p0_rdat_1129 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1130 = {_zz_shareBuffer_sbuf_p0_rdat_1131,_zz_shareBuffer_sbuf_p0_rdat_1132};
  assign _zz_shareBuffer_sbuf_p0_rdat_1242 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1243 = {_zz_shareBuffer_sbuf_p0_rdat_1244,_zz_shareBuffer_sbuf_p0_rdat_1245};
  assign _zz_shareBuffer_sbuf_p0_rdat_1355 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1356 = {_zz_shareBuffer_sbuf_p0_rdat_1357,_zz_shareBuffer_sbuf_p0_rdat_1358};
  assign _zz_shareBuffer_sbuf_p0_rdat_1467 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1468 = {_zz_shareBuffer_sbuf_p0_rdat_1469,_zz_shareBuffer_sbuf_p0_rdat_1470};
  assign _zz_shareBuffer_sbuf_p0_rdat_1579 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1580 = {_zz_shareBuffer_sbuf_p0_rdat_1581,_zz_shareBuffer_sbuf_p0_rdat_1582};
  assign _zz_shareBuffer_sbuf_p0_rdat_1689 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1690 = {_zz_shareBuffer_sbuf_p0_rdat_1691,_zz_shareBuffer_sbuf_p0_rdat_1692};
  assign _zz_shareBuffer_sbuf_p0_rdat_6 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_7 = {_zz_shareBuffer_sbuf_p0_rdat_8,_zz_shareBuffer_sbuf_p0_rdat_9};
  assign _zz_shareBuffer_sbuf_p0_rdat_115 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_116 = {_zz_shareBuffer_sbuf_p0_rdat_117,_zz_shareBuffer_sbuf_p0_rdat_118};
  assign _zz_shareBuffer_sbuf_p0_rdat_226 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_227 = {_zz_shareBuffer_sbuf_p0_rdat_228,_zz_shareBuffer_sbuf_p0_rdat_229};
  assign _zz_shareBuffer_sbuf_p0_rdat_337 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_338 = {_zz_shareBuffer_sbuf_p0_rdat_339,_zz_shareBuffer_sbuf_p0_rdat_340};
  assign _zz_shareBuffer_sbuf_p0_rdat_450 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_451 = {_zz_shareBuffer_sbuf_p0_rdat_452,_zz_shareBuffer_sbuf_p0_rdat_453};
  assign _zz_shareBuffer_sbuf_p0_rdat_563 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_564 = {_zz_shareBuffer_sbuf_p0_rdat_565,_zz_shareBuffer_sbuf_p0_rdat_566};
  assign _zz_shareBuffer_sbuf_p0_rdat_676 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_677 = {_zz_shareBuffer_sbuf_p0_rdat_678,_zz_shareBuffer_sbuf_p0_rdat_679};
  assign _zz_shareBuffer_sbuf_p0_rdat_789 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_790 = {_zz_shareBuffer_sbuf_p0_rdat_791,_zz_shareBuffer_sbuf_p0_rdat_792};
  assign _zz_shareBuffer_sbuf_p0_rdat_904 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_905 = {_zz_shareBuffer_sbuf_p0_rdat_906,_zz_shareBuffer_sbuf_p0_rdat_907};
  assign _zz_shareBuffer_sbuf_p0_rdat_1017 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1018 = {_zz_shareBuffer_sbuf_p0_rdat_1019,_zz_shareBuffer_sbuf_p0_rdat_1020};
  assign _zz_shareBuffer_sbuf_p0_rdat_1131 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1132 = {_zz_shareBuffer_sbuf_p0_rdat_1133,_zz_shareBuffer_sbuf_p0_rdat_1134};
  assign _zz_shareBuffer_sbuf_p0_rdat_1244 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1245 = {_zz_shareBuffer_sbuf_p0_rdat_1246,_zz_shareBuffer_sbuf_p0_rdat_1247};
  assign _zz_shareBuffer_sbuf_p0_rdat_1357 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1358 = {_zz_shareBuffer_sbuf_p0_rdat_1359,_zz_shareBuffer_sbuf_p0_rdat_1360};
  assign _zz_shareBuffer_sbuf_p0_rdat_1469 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1470 = {_zz_shareBuffer_sbuf_p0_rdat_1471,_zz_shareBuffer_sbuf_p0_rdat_1472};
  assign _zz_shareBuffer_sbuf_p0_rdat_1581 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1582 = {_zz_shareBuffer_sbuf_p0_rdat_1583,_zz_shareBuffer_sbuf_p0_rdat_1584};
  assign _zz_shareBuffer_sbuf_p0_rdat_1691 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1692 = {_zz_shareBuffer_sbuf_p0_rdat_1693,_zz_shareBuffer_sbuf_p0_rdat_1694};
  assign _zz_shareBuffer_sbuf_p0_rdat_8 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_9 = {_zz_shareBuffer_sbuf_p0_rdat_10,_zz_shareBuffer_sbuf_p0_rdat_11};
  assign _zz_shareBuffer_sbuf_p0_rdat_117 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_118 = {_zz_shareBuffer_sbuf_p0_rdat_119,_zz_shareBuffer_sbuf_p0_rdat_120};
  assign _zz_shareBuffer_sbuf_p0_rdat_228 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_229 = {_zz_shareBuffer_sbuf_p0_rdat_230,_zz_shareBuffer_sbuf_p0_rdat_231};
  assign _zz_shareBuffer_sbuf_p0_rdat_339 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_340 = {_zz_shareBuffer_sbuf_p0_rdat_341,_zz_shareBuffer_sbuf_p0_rdat_342};
  assign _zz_shareBuffer_sbuf_p0_rdat_452 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_453 = {_zz_shareBuffer_sbuf_p0_rdat_454,_zz_shareBuffer_sbuf_p0_rdat_455};
  assign _zz_shareBuffer_sbuf_p0_rdat_565 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_566 = {_zz_shareBuffer_sbuf_p0_rdat_567,_zz_shareBuffer_sbuf_p0_rdat_568};
  assign _zz_shareBuffer_sbuf_p0_rdat_678 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_679 = {_zz_shareBuffer_sbuf_p0_rdat_680,_zz_shareBuffer_sbuf_p0_rdat_681};
  assign _zz_shareBuffer_sbuf_p0_rdat_791 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_792 = {_zz_shareBuffer_sbuf_p0_rdat_793,_zz_shareBuffer_sbuf_p0_rdat_794};
  assign _zz_shareBuffer_sbuf_p0_rdat_906 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_907 = {_zz_shareBuffer_sbuf_p0_rdat_908,_zz_shareBuffer_sbuf_p0_rdat_909};
  assign _zz_shareBuffer_sbuf_p0_rdat_1019 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1020 = {_zz_shareBuffer_sbuf_p0_rdat_1021,_zz_shareBuffer_sbuf_p0_rdat_1022};
  assign _zz_shareBuffer_sbuf_p0_rdat_1133 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1134 = {_zz_shareBuffer_sbuf_p0_rdat_1135,_zz_shareBuffer_sbuf_p0_rdat_1136};
  assign _zz_shareBuffer_sbuf_p0_rdat_1246 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1247 = {_zz_shareBuffer_sbuf_p0_rdat_1248,_zz_shareBuffer_sbuf_p0_rdat_1249};
  assign _zz_shareBuffer_sbuf_p0_rdat_1359 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1360 = {_zz_shareBuffer_sbuf_p0_rdat_1361,_zz_shareBuffer_sbuf_p0_rdat_1362};
  assign _zz_shareBuffer_sbuf_p0_rdat_1471 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1472 = {_zz_shareBuffer_sbuf_p0_rdat_1473,_zz_shareBuffer_sbuf_p0_rdat_1474};
  assign _zz_shareBuffer_sbuf_p0_rdat_1583 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1584 = {_zz_shareBuffer_sbuf_p0_rdat_1585,_zz_shareBuffer_sbuf_p0_rdat_1586};
  assign _zz_shareBuffer_sbuf_p0_rdat_1693 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1694 = {_zz_shareBuffer_sbuf_p0_rdat_1695,_zz_shareBuffer_sbuf_p0_rdat_1696};
  assign _zz_shareBuffer_sbuf_p0_rdat_10 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_11 = {_zz_shareBuffer_sbuf_p0_rdat_12,_zz_shareBuffer_sbuf_p0_rdat_13};
  assign _zz_shareBuffer_sbuf_p0_rdat_119 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_120 = {_zz_shareBuffer_sbuf_p0_rdat_121,_zz_shareBuffer_sbuf_p0_rdat_122};
  assign _zz_shareBuffer_sbuf_p0_rdat_230 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_231 = {_zz_shareBuffer_sbuf_p0_rdat_232,_zz_shareBuffer_sbuf_p0_rdat_233};
  assign _zz_shareBuffer_sbuf_p0_rdat_341 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_342 = {_zz_shareBuffer_sbuf_p0_rdat_343,_zz_shareBuffer_sbuf_p0_rdat_344};
  assign _zz_shareBuffer_sbuf_p0_rdat_454 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_455 = {_zz_shareBuffer_sbuf_p0_rdat_456,_zz_shareBuffer_sbuf_p0_rdat_457};
  assign _zz_shareBuffer_sbuf_p0_rdat_567 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_568 = {_zz_shareBuffer_sbuf_p0_rdat_569,_zz_shareBuffer_sbuf_p0_rdat_570};
  assign _zz_shareBuffer_sbuf_p0_rdat_680 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_681 = {_zz_shareBuffer_sbuf_p0_rdat_682,_zz_shareBuffer_sbuf_p0_rdat_683};
  assign _zz_shareBuffer_sbuf_p0_rdat_793 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_794 = {_zz_shareBuffer_sbuf_p0_rdat_795,_zz_shareBuffer_sbuf_p0_rdat_796};
  assign _zz_shareBuffer_sbuf_p0_rdat_908 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_909 = {_zz_shareBuffer_sbuf_p0_rdat_910,_zz_shareBuffer_sbuf_p0_rdat_911};
  assign _zz_shareBuffer_sbuf_p0_rdat_1021 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1022 = {_zz_shareBuffer_sbuf_p0_rdat_1023,_zz_shareBuffer_sbuf_p0_rdat_1024};
  assign _zz_shareBuffer_sbuf_p0_rdat_1135 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1136 = {_zz_shareBuffer_sbuf_p0_rdat_1137,_zz_shareBuffer_sbuf_p0_rdat_1138};
  assign _zz_shareBuffer_sbuf_p0_rdat_1248 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1249 = {_zz_shareBuffer_sbuf_p0_rdat_1250,_zz_shareBuffer_sbuf_p0_rdat_1251};
  assign _zz_shareBuffer_sbuf_p0_rdat_1361 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1362 = {_zz_shareBuffer_sbuf_p0_rdat_1363,_zz_shareBuffer_sbuf_p0_rdat_1364};
  assign _zz_shareBuffer_sbuf_p0_rdat_1473 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1474 = {_zz_shareBuffer_sbuf_p0_rdat_1475,_zz_shareBuffer_sbuf_p0_rdat_1476};
  assign _zz_shareBuffer_sbuf_p0_rdat_1585 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1586 = {_zz_shareBuffer_sbuf_p0_rdat_1587,_zz_shareBuffer_sbuf_p0_rdat_1588};
  assign _zz_shareBuffer_sbuf_p0_rdat_1695 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1696 = {_zz_shareBuffer_sbuf_p0_rdat_1697,_zz_shareBuffer_sbuf_p0_rdat_1698};
  assign _zz_shareBuffer_sbuf_p0_rdat_12 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_13 = {_zz_shareBuffer_sbuf_p0_rdat_14,_zz_shareBuffer_sbuf_p0_rdat_15};
  assign _zz_shareBuffer_sbuf_p0_rdat_121 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_122 = {_zz_shareBuffer_sbuf_p0_rdat_123,_zz_shareBuffer_sbuf_p0_rdat_124};
  assign _zz_shareBuffer_sbuf_p0_rdat_232 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_233 = {_zz_shareBuffer_sbuf_p0_rdat_234,_zz_shareBuffer_sbuf_p0_rdat_235};
  assign _zz_shareBuffer_sbuf_p0_rdat_343 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_344 = {_zz_shareBuffer_sbuf_p0_rdat_345,_zz_shareBuffer_sbuf_p0_rdat_346};
  assign _zz_shareBuffer_sbuf_p0_rdat_456 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_457 = {_zz_shareBuffer_sbuf_p0_rdat_458,_zz_shareBuffer_sbuf_p0_rdat_459};
  assign _zz_shareBuffer_sbuf_p0_rdat_569 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_570 = {_zz_shareBuffer_sbuf_p0_rdat_571,_zz_shareBuffer_sbuf_p0_rdat_572};
  assign _zz_shareBuffer_sbuf_p0_rdat_682 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_683 = {_zz_shareBuffer_sbuf_p0_rdat_684,_zz_shareBuffer_sbuf_p0_rdat_685};
  assign _zz_shareBuffer_sbuf_p0_rdat_795 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_796 = {_zz_shareBuffer_sbuf_p0_rdat_797,_zz_shareBuffer_sbuf_p0_rdat_798};
  assign _zz_shareBuffer_sbuf_p0_rdat_910 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_911 = {_zz_shareBuffer_sbuf_p0_rdat_912,_zz_shareBuffer_sbuf_p0_rdat_913};
  assign _zz_shareBuffer_sbuf_p0_rdat_1023 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1024 = {_zz_shareBuffer_sbuf_p0_rdat_1025,_zz_shareBuffer_sbuf_p0_rdat_1026};
  assign _zz_shareBuffer_sbuf_p0_rdat_1137 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1138 = {_zz_shareBuffer_sbuf_p0_rdat_1139,_zz_shareBuffer_sbuf_p0_rdat_1140};
  assign _zz_shareBuffer_sbuf_p0_rdat_1250 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1251 = {_zz_shareBuffer_sbuf_p0_rdat_1252,_zz_shareBuffer_sbuf_p0_rdat_1253};
  assign _zz_shareBuffer_sbuf_p0_rdat_1363 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1364 = {_zz_shareBuffer_sbuf_p0_rdat_1365,_zz_shareBuffer_sbuf_p0_rdat_1366};
  assign _zz_shareBuffer_sbuf_p0_rdat_1475 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1476 = {_zz_shareBuffer_sbuf_p0_rdat_1477,_zz_shareBuffer_sbuf_p0_rdat_1478};
  assign _zz_shareBuffer_sbuf_p0_rdat_1587 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1588 = {_zz_shareBuffer_sbuf_p0_rdat_1589,_zz_shareBuffer_sbuf_p0_rdat_1590};
  assign _zz_shareBuffer_sbuf_p0_rdat_1697 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1698 = {_zz_shareBuffer_sbuf_p0_rdat_1699,_zz_shareBuffer_sbuf_p0_rdat_1700};
  assign _zz_shareBuffer_sbuf_p0_rdat_14 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_15 = {_zz_shareBuffer_sbuf_p0_rdat_16,_zz_shareBuffer_sbuf_p0_rdat_17};
  assign _zz_shareBuffer_sbuf_p0_rdat_123 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_124 = {_zz_shareBuffer_sbuf_p0_rdat_125,_zz_shareBuffer_sbuf_p0_rdat_126};
  assign _zz_shareBuffer_sbuf_p0_rdat_234 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_235 = {_zz_shareBuffer_sbuf_p0_rdat_236,_zz_shareBuffer_sbuf_p0_rdat_237};
  assign _zz_shareBuffer_sbuf_p0_rdat_345 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_346 = {_zz_shareBuffer_sbuf_p0_rdat_347,_zz_shareBuffer_sbuf_p0_rdat_348};
  assign _zz_shareBuffer_sbuf_p0_rdat_458 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_459 = {_zz_shareBuffer_sbuf_p0_rdat_460,_zz_shareBuffer_sbuf_p0_rdat_461};
  assign _zz_shareBuffer_sbuf_p0_rdat_571 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_572 = {_zz_shareBuffer_sbuf_p0_rdat_573,_zz_shareBuffer_sbuf_p0_rdat_574};
  assign _zz_shareBuffer_sbuf_p0_rdat_684 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_685 = {_zz_shareBuffer_sbuf_p0_rdat_686,_zz_shareBuffer_sbuf_p0_rdat_687};
  assign _zz_shareBuffer_sbuf_p0_rdat_797 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_798 = {_zz_shareBuffer_sbuf_p0_rdat_799,_zz_shareBuffer_sbuf_p0_rdat_800};
  assign _zz_shareBuffer_sbuf_p0_rdat_912 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_913 = {_zz_shareBuffer_sbuf_p0_rdat_914,_zz_shareBuffer_sbuf_p0_rdat_915};
  assign _zz_shareBuffer_sbuf_p0_rdat_1025 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1026 = {_zz_shareBuffer_sbuf_p0_rdat_1027,_zz_shareBuffer_sbuf_p0_rdat_1028};
  assign _zz_shareBuffer_sbuf_p0_rdat_1139 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1140 = {_zz_shareBuffer_sbuf_p0_rdat_1141,_zz_shareBuffer_sbuf_p0_rdat_1142};
  assign _zz_shareBuffer_sbuf_p0_rdat_1252 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1253 = {_zz_shareBuffer_sbuf_p0_rdat_1254,_zz_shareBuffer_sbuf_p0_rdat_1255};
  assign _zz_shareBuffer_sbuf_p0_rdat_1365 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1366 = {_zz_shareBuffer_sbuf_p0_rdat_1367,_zz_shareBuffer_sbuf_p0_rdat_1368};
  assign _zz_shareBuffer_sbuf_p0_rdat_1477 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1478 = {_zz_shareBuffer_sbuf_p0_rdat_1479,_zz_shareBuffer_sbuf_p0_rdat_1480};
  assign _zz_shareBuffer_sbuf_p0_rdat_1589 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1590 = {_zz_shareBuffer_sbuf_p0_rdat_1591,_zz_shareBuffer_sbuf_p0_rdat_1592};
  assign _zz_shareBuffer_sbuf_p0_rdat_1699 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1700 = {_zz_shareBuffer_sbuf_p0_rdat_1701,_zz_shareBuffer_sbuf_p0_rdat_1702};
  assign _zz_shareBuffer_sbuf_p0_rdat_16 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_17 = {_zz_shareBuffer_sbuf_p0_rdat_18,_zz_shareBuffer_sbuf_p0_rdat_19};
  assign _zz_shareBuffer_sbuf_p0_rdat_125 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_126 = {_zz_shareBuffer_sbuf_p0_rdat_127,_zz_shareBuffer_sbuf_p0_rdat_128};
  assign _zz_shareBuffer_sbuf_p0_rdat_236 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_237 = {_zz_shareBuffer_sbuf_p0_rdat_238,_zz_shareBuffer_sbuf_p0_rdat_239};
  assign _zz_shareBuffer_sbuf_p0_rdat_347 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_348 = {_zz_shareBuffer_sbuf_p0_rdat_349,_zz_shareBuffer_sbuf_p0_rdat_350};
  assign _zz_shareBuffer_sbuf_p0_rdat_460 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_461 = {_zz_shareBuffer_sbuf_p0_rdat_462,_zz_shareBuffer_sbuf_p0_rdat_463};
  assign _zz_shareBuffer_sbuf_p0_rdat_573 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_574 = {_zz_shareBuffer_sbuf_p0_rdat_575,_zz_shareBuffer_sbuf_p0_rdat_576};
  assign _zz_shareBuffer_sbuf_p0_rdat_686 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_687 = {_zz_shareBuffer_sbuf_p0_rdat_688,_zz_shareBuffer_sbuf_p0_rdat_689};
  assign _zz_shareBuffer_sbuf_p0_rdat_799 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_800 = {_zz_shareBuffer_sbuf_p0_rdat_801,_zz_shareBuffer_sbuf_p0_rdat_802};
  assign _zz_shareBuffer_sbuf_p0_rdat_914 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_915 = {_zz_shareBuffer_sbuf_p0_rdat_916,_zz_shareBuffer_sbuf_p0_rdat_917};
  assign _zz_shareBuffer_sbuf_p0_rdat_1027 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1028 = {_zz_shareBuffer_sbuf_p0_rdat_1029,_zz_shareBuffer_sbuf_p0_rdat_1030};
  assign _zz_shareBuffer_sbuf_p0_rdat_1141 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1142 = {_zz_shareBuffer_sbuf_p0_rdat_1143,_zz_shareBuffer_sbuf_p0_rdat_1144};
  assign _zz_shareBuffer_sbuf_p0_rdat_1254 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1255 = {_zz_shareBuffer_sbuf_p0_rdat_1256,_zz_shareBuffer_sbuf_p0_rdat_1257};
  assign _zz_shareBuffer_sbuf_p0_rdat_1367 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1368 = {_zz_shareBuffer_sbuf_p0_rdat_1369,_zz_shareBuffer_sbuf_p0_rdat_1370};
  assign _zz_shareBuffer_sbuf_p0_rdat_1479 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1480 = {_zz_shareBuffer_sbuf_p0_rdat_1481,_zz_shareBuffer_sbuf_p0_rdat_1482};
  assign _zz_shareBuffer_sbuf_p0_rdat_1591 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1592 = {_zz_shareBuffer_sbuf_p0_rdat_1593,_zz_shareBuffer_sbuf_p0_rdat_1594};
  assign _zz_shareBuffer_sbuf_p0_rdat_1701 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1702 = {_zz_shareBuffer_sbuf_p0_rdat_1703,_zz_shareBuffer_sbuf_p0_rdat_1704};
  assign _zz_shareBuffer_sbuf_p0_rdat_18 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_19 = {_zz_shareBuffer_sbuf_p0_rdat_20,_zz_shareBuffer_sbuf_p0_rdat_21};
  assign _zz_shareBuffer_sbuf_p0_rdat_127 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_128 = {_zz_shareBuffer_sbuf_p0_rdat_129,_zz_shareBuffer_sbuf_p0_rdat_130};
  assign _zz_shareBuffer_sbuf_p0_rdat_238 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_239 = {_zz_shareBuffer_sbuf_p0_rdat_240,_zz_shareBuffer_sbuf_p0_rdat_241};
  assign _zz_shareBuffer_sbuf_p0_rdat_349 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_350 = {_zz_shareBuffer_sbuf_p0_rdat_351,_zz_shareBuffer_sbuf_p0_rdat_352};
  assign _zz_shareBuffer_sbuf_p0_rdat_462 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_463 = {_zz_shareBuffer_sbuf_p0_rdat_464,_zz_shareBuffer_sbuf_p0_rdat_465};
  assign _zz_shareBuffer_sbuf_p0_rdat_575 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_576 = {_zz_shareBuffer_sbuf_p0_rdat_577,_zz_shareBuffer_sbuf_p0_rdat_578};
  assign _zz_shareBuffer_sbuf_p0_rdat_688 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_689 = {_zz_shareBuffer_sbuf_p0_rdat_690,_zz_shareBuffer_sbuf_p0_rdat_691};
  assign _zz_shareBuffer_sbuf_p0_rdat_801 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_802 = {_zz_shareBuffer_sbuf_p0_rdat_803,_zz_shareBuffer_sbuf_p0_rdat_804};
  assign _zz_shareBuffer_sbuf_p0_rdat_916 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_917 = {_zz_shareBuffer_sbuf_p0_rdat_918,_zz_shareBuffer_sbuf_p0_rdat_919};
  assign _zz_shareBuffer_sbuf_p0_rdat_1029 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1030 = {_zz_shareBuffer_sbuf_p0_rdat_1031,_zz_shareBuffer_sbuf_p0_rdat_1032};
  assign _zz_shareBuffer_sbuf_p0_rdat_1143 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1144 = {_zz_shareBuffer_sbuf_p0_rdat_1145,_zz_shareBuffer_sbuf_p0_rdat_1146};
  assign _zz_shareBuffer_sbuf_p0_rdat_1256 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1257 = {_zz_shareBuffer_sbuf_p0_rdat_1258,_zz_shareBuffer_sbuf_p0_rdat_1259};
  assign _zz_shareBuffer_sbuf_p0_rdat_1369 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1370 = {_zz_shareBuffer_sbuf_p0_rdat_1371,_zz_shareBuffer_sbuf_p0_rdat_1372};
  assign _zz_shareBuffer_sbuf_p0_rdat_1481 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1482 = {_zz_shareBuffer_sbuf_p0_rdat_1483,_zz_shareBuffer_sbuf_p0_rdat_1484};
  assign _zz_shareBuffer_sbuf_p0_rdat_1593 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1594 = {_zz_shareBuffer_sbuf_p0_rdat_1595,_zz_shareBuffer_sbuf_p0_rdat_1596};
  assign _zz_shareBuffer_sbuf_p0_rdat_1703 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1704 = {_zz_shareBuffer_sbuf_p0_rdat_1705,_zz_shareBuffer_sbuf_p0_rdat_1706};
  assign _zz_shareBuffer_sbuf_p0_rdat_20 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_21 = {_zz_shareBuffer_sbuf_p0_rdat_22,_zz_shareBuffer_sbuf_p0_rdat_23};
  assign _zz_shareBuffer_sbuf_p0_rdat_129 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_130 = {_zz_shareBuffer_sbuf_p0_rdat_131,_zz_shareBuffer_sbuf_p0_rdat_132};
  assign _zz_shareBuffer_sbuf_p0_rdat_240 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_241 = {_zz_shareBuffer_sbuf_p0_rdat_242,_zz_shareBuffer_sbuf_p0_rdat_243};
  assign _zz_shareBuffer_sbuf_p0_rdat_351 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_352 = {_zz_shareBuffer_sbuf_p0_rdat_353,_zz_shareBuffer_sbuf_p0_rdat_354};
  assign _zz_shareBuffer_sbuf_p0_rdat_464 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_465 = {_zz_shareBuffer_sbuf_p0_rdat_466,_zz_shareBuffer_sbuf_p0_rdat_467};
  assign _zz_shareBuffer_sbuf_p0_rdat_577 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_578 = {_zz_shareBuffer_sbuf_p0_rdat_579,_zz_shareBuffer_sbuf_p0_rdat_580};
  assign _zz_shareBuffer_sbuf_p0_rdat_690 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_691 = {_zz_shareBuffer_sbuf_p0_rdat_692,_zz_shareBuffer_sbuf_p0_rdat_693};
  assign _zz_shareBuffer_sbuf_p0_rdat_803 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_804 = {_zz_shareBuffer_sbuf_p0_rdat_805,_zz_shareBuffer_sbuf_p0_rdat_806};
  assign _zz_shareBuffer_sbuf_p0_rdat_918 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_919 = {_zz_shareBuffer_sbuf_p0_rdat_920,_zz_shareBuffer_sbuf_p0_rdat_921};
  assign _zz_shareBuffer_sbuf_p0_rdat_1031 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1032 = {_zz_shareBuffer_sbuf_p0_rdat_1033,_zz_shareBuffer_sbuf_p0_rdat_1034};
  assign _zz_shareBuffer_sbuf_p0_rdat_1145 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1146 = {_zz_shareBuffer_sbuf_p0_rdat_1147,_zz_shareBuffer_sbuf_p0_rdat_1148};
  assign _zz_shareBuffer_sbuf_p0_rdat_1258 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1259 = {_zz_shareBuffer_sbuf_p0_rdat_1260,_zz_shareBuffer_sbuf_p0_rdat_1261};
  assign _zz_shareBuffer_sbuf_p0_rdat_1371 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1372 = {_zz_shareBuffer_sbuf_p0_rdat_1373,_zz_shareBuffer_sbuf_p0_rdat_1374};
  assign _zz_shareBuffer_sbuf_p0_rdat_1483 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1484 = {_zz_shareBuffer_sbuf_p0_rdat_1485,_zz_shareBuffer_sbuf_p0_rdat_1486};
  assign _zz_shareBuffer_sbuf_p0_rdat_1595 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1596 = {_zz_shareBuffer_sbuf_p0_rdat_1597,_zz_shareBuffer_sbuf_p0_rdat_1598};
  assign _zz_shareBuffer_sbuf_p0_rdat_1705 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1706 = {_zz_shareBuffer_sbuf_p0_rdat_1707,_zz_shareBuffer_sbuf_p0_rdat_1708};
  assign _zz_shareBuffer_sbuf_p0_rdat_22 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_23 = {_zz_shareBuffer_sbuf_p0_rdat_24,_zz_shareBuffer_sbuf_p0_rdat_25};
  assign _zz_shareBuffer_sbuf_p0_rdat_131 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_132 = {_zz_shareBuffer_sbuf_p0_rdat_133,_zz_shareBuffer_sbuf_p0_rdat_134};
  assign _zz_shareBuffer_sbuf_p0_rdat_242 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_243 = {_zz_shareBuffer_sbuf_p0_rdat_244,_zz_shareBuffer_sbuf_p0_rdat_245};
  assign _zz_shareBuffer_sbuf_p0_rdat_353 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_354 = {_zz_shareBuffer_sbuf_p0_rdat_355,_zz_shareBuffer_sbuf_p0_rdat_356};
  assign _zz_shareBuffer_sbuf_p0_rdat_466 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_467 = {_zz_shareBuffer_sbuf_p0_rdat_468,_zz_shareBuffer_sbuf_p0_rdat_469};
  assign _zz_shareBuffer_sbuf_p0_rdat_579 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_580 = {_zz_shareBuffer_sbuf_p0_rdat_581,_zz_shareBuffer_sbuf_p0_rdat_582};
  assign _zz_shareBuffer_sbuf_p0_rdat_692 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_693 = {_zz_shareBuffer_sbuf_p0_rdat_694,_zz_shareBuffer_sbuf_p0_rdat_695};
  assign _zz_shareBuffer_sbuf_p0_rdat_805 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_806 = {_zz_shareBuffer_sbuf_p0_rdat_807,_zz_shareBuffer_sbuf_p0_rdat_808};
  assign _zz_shareBuffer_sbuf_p0_rdat_920 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_921 = {_zz_shareBuffer_sbuf_p0_rdat_922,_zz_shareBuffer_sbuf_p0_rdat_923};
  assign _zz_shareBuffer_sbuf_p0_rdat_1033 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1034 = {_zz_shareBuffer_sbuf_p0_rdat_1035,_zz_shareBuffer_sbuf_p0_rdat_1036};
  assign _zz_shareBuffer_sbuf_p0_rdat_1147 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1148 = {_zz_shareBuffer_sbuf_p0_rdat_1149,_zz_shareBuffer_sbuf_p0_rdat_1150};
  assign _zz_shareBuffer_sbuf_p0_rdat_1260 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1261 = {_zz_shareBuffer_sbuf_p0_rdat_1262,_zz_shareBuffer_sbuf_p0_rdat_1263};
  assign _zz_shareBuffer_sbuf_p0_rdat_1373 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1374 = {_zz_shareBuffer_sbuf_p0_rdat_1375,_zz_shareBuffer_sbuf_p0_rdat_1376};
  assign _zz_shareBuffer_sbuf_p0_rdat_1485 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1486 = {_zz_shareBuffer_sbuf_p0_rdat_1487,_zz_shareBuffer_sbuf_p0_rdat_1488};
  assign _zz_shareBuffer_sbuf_p0_rdat_1597 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1598 = {_zz_shareBuffer_sbuf_p0_rdat_1599,_zz_shareBuffer_sbuf_p0_rdat_1600};
  assign _zz_shareBuffer_sbuf_p0_rdat_1707 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1708 = {_zz_shareBuffer_sbuf_p0_rdat_1709,_zz_shareBuffer_sbuf_p0_rdat_1710};
  assign _zz_shareBuffer_sbuf_p0_rdat_24 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_25 = {_zz_shareBuffer_sbuf_p0_rdat_26,_zz_shareBuffer_sbuf_p0_rdat_27};
  assign _zz_shareBuffer_sbuf_p0_rdat_133 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_134 = {_zz_shareBuffer_sbuf_p0_rdat_135,_zz_shareBuffer_sbuf_p0_rdat_136};
  assign _zz_shareBuffer_sbuf_p0_rdat_244 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_245 = {_zz_shareBuffer_sbuf_p0_rdat_246,_zz_shareBuffer_sbuf_p0_rdat_247};
  assign _zz_shareBuffer_sbuf_p0_rdat_355 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_356 = {_zz_shareBuffer_sbuf_p0_rdat_357,_zz_shareBuffer_sbuf_p0_rdat_358};
  assign _zz_shareBuffer_sbuf_p0_rdat_468 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_469 = {_zz_shareBuffer_sbuf_p0_rdat_470,_zz_shareBuffer_sbuf_p0_rdat_471};
  assign _zz_shareBuffer_sbuf_p0_rdat_581 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_582 = {_zz_shareBuffer_sbuf_p0_rdat_583,_zz_shareBuffer_sbuf_p0_rdat_584};
  assign _zz_shareBuffer_sbuf_p0_rdat_694 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_695 = {_zz_shareBuffer_sbuf_p0_rdat_696,_zz_shareBuffer_sbuf_p0_rdat_697};
  assign _zz_shareBuffer_sbuf_p0_rdat_807 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_808 = {_zz_shareBuffer_sbuf_p0_rdat_809,_zz_shareBuffer_sbuf_p0_rdat_810};
  assign _zz_shareBuffer_sbuf_p0_rdat_922 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_923 = {_zz_shareBuffer_sbuf_p0_rdat_924,_zz_shareBuffer_sbuf_p0_rdat_925};
  assign _zz_shareBuffer_sbuf_p0_rdat_1035 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1036 = {_zz_shareBuffer_sbuf_p0_rdat_1037,_zz_shareBuffer_sbuf_p0_rdat_1038};
  assign _zz_shareBuffer_sbuf_p0_rdat_1149 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1150 = {_zz_shareBuffer_sbuf_p0_rdat_1151,_zz_shareBuffer_sbuf_p0_rdat_1152};
  assign _zz_shareBuffer_sbuf_p0_rdat_1262 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1263 = {_zz_shareBuffer_sbuf_p0_rdat_1264,_zz_shareBuffer_sbuf_p0_rdat_1265};
  assign _zz_shareBuffer_sbuf_p0_rdat_1375 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1376 = {_zz_shareBuffer_sbuf_p0_rdat_1377,_zz_shareBuffer_sbuf_p0_rdat_1378};
  assign _zz_shareBuffer_sbuf_p0_rdat_1487 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1488 = {_zz_shareBuffer_sbuf_p0_rdat_1489,_zz_shareBuffer_sbuf_p0_rdat_1490};
  assign _zz_shareBuffer_sbuf_p0_rdat_1599 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1600 = {_zz_shareBuffer_sbuf_p0_rdat_1601,_zz_shareBuffer_sbuf_p0_rdat_1602};
  assign _zz_shareBuffer_sbuf_p0_rdat_1709 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1710 = {_zz_shareBuffer_sbuf_p0_rdat_1711,_zz_shareBuffer_sbuf_p0_rdat_1712};
  assign _zz_shareBuffer_sbuf_p0_rdat_26 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_27 = {_zz_shareBuffer_sbuf_p0_rdat_28,_zz_shareBuffer_sbuf_p0_rdat_29};
  assign _zz_shareBuffer_sbuf_p0_rdat_135 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_136 = {_zz_shareBuffer_sbuf_p0_rdat_137,_zz_shareBuffer_sbuf_p0_rdat_138};
  assign _zz_shareBuffer_sbuf_p0_rdat_246 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_247 = {_zz_shareBuffer_sbuf_p0_rdat_248,_zz_shareBuffer_sbuf_p0_rdat_249};
  assign _zz_shareBuffer_sbuf_p0_rdat_357 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_358 = {_zz_shareBuffer_sbuf_p0_rdat_359,_zz_shareBuffer_sbuf_p0_rdat_360};
  assign _zz_shareBuffer_sbuf_p0_rdat_470 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_471 = {_zz_shareBuffer_sbuf_p0_rdat_472,_zz_shareBuffer_sbuf_p0_rdat_473};
  assign _zz_shareBuffer_sbuf_p0_rdat_583 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_584 = {_zz_shareBuffer_sbuf_p0_rdat_585,_zz_shareBuffer_sbuf_p0_rdat_586};
  assign _zz_shareBuffer_sbuf_p0_rdat_696 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_697 = {_zz_shareBuffer_sbuf_p0_rdat_698,_zz_shareBuffer_sbuf_p0_rdat_699};
  assign _zz_shareBuffer_sbuf_p0_rdat_809 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_810 = {_zz_shareBuffer_sbuf_p0_rdat_811,_zz_shareBuffer_sbuf_p0_rdat_812};
  assign _zz_shareBuffer_sbuf_p0_rdat_924 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_925 = {_zz_shareBuffer_sbuf_p0_rdat_926,_zz_shareBuffer_sbuf_p0_rdat_927};
  assign _zz_shareBuffer_sbuf_p0_rdat_1037 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1038 = {_zz_shareBuffer_sbuf_p0_rdat_1039,_zz_shareBuffer_sbuf_p0_rdat_1040};
  assign _zz_shareBuffer_sbuf_p0_rdat_1151 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1152 = {_zz_shareBuffer_sbuf_p0_rdat_1153,_zz_shareBuffer_sbuf_p0_rdat_1154};
  assign _zz_shareBuffer_sbuf_p0_rdat_1264 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1265 = {_zz_shareBuffer_sbuf_p0_rdat_1266,_zz_shareBuffer_sbuf_p0_rdat_1267};
  assign _zz_shareBuffer_sbuf_p0_rdat_1377 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1378 = {_zz_shareBuffer_sbuf_p0_rdat_1379,_zz_shareBuffer_sbuf_p0_rdat_1380};
  assign _zz_shareBuffer_sbuf_p0_rdat_1489 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1490 = {_zz_shareBuffer_sbuf_p0_rdat_1491,_zz_shareBuffer_sbuf_p0_rdat_1492};
  assign _zz_shareBuffer_sbuf_p0_rdat_1601 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1602 = {_zz_shareBuffer_sbuf_p0_rdat_1603,_zz_shareBuffer_sbuf_p0_rdat_1604};
  assign _zz_shareBuffer_sbuf_p0_rdat_1711 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1712 = {_zz_shareBuffer_sbuf_p0_rdat_1713,_zz_shareBuffer_sbuf_p0_rdat_1714};
  assign _zz_shareBuffer_sbuf_p0_rdat_28 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_29 = {_zz_shareBuffer_sbuf_p0_rdat_30,_zz_shareBuffer_sbuf_p0_rdat_31};
  assign _zz_shareBuffer_sbuf_p0_rdat_137 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_138 = {_zz_shareBuffer_sbuf_p0_rdat_139,_zz_shareBuffer_sbuf_p0_rdat_140};
  assign _zz_shareBuffer_sbuf_p0_rdat_248 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_249 = {_zz_shareBuffer_sbuf_p0_rdat_250,_zz_shareBuffer_sbuf_p0_rdat_251};
  assign _zz_shareBuffer_sbuf_p0_rdat_359 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_360 = {_zz_shareBuffer_sbuf_p0_rdat_361,_zz_shareBuffer_sbuf_p0_rdat_362};
  assign _zz_shareBuffer_sbuf_p0_rdat_472 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_473 = {_zz_shareBuffer_sbuf_p0_rdat_474,_zz_shareBuffer_sbuf_p0_rdat_475};
  assign _zz_shareBuffer_sbuf_p0_rdat_585 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_586 = {_zz_shareBuffer_sbuf_p0_rdat_587,_zz_shareBuffer_sbuf_p0_rdat_588};
  assign _zz_shareBuffer_sbuf_p0_rdat_698 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_699 = {_zz_shareBuffer_sbuf_p0_rdat_700,_zz_shareBuffer_sbuf_p0_rdat_701};
  assign _zz_shareBuffer_sbuf_p0_rdat_811 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_812 = {_zz_shareBuffer_sbuf_p0_rdat_813,_zz_shareBuffer_sbuf_p0_rdat_814};
  assign _zz_shareBuffer_sbuf_p0_rdat_926 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_927 = {_zz_shareBuffer_sbuf_p0_rdat_928,_zz_shareBuffer_sbuf_p0_rdat_929};
  assign _zz_shareBuffer_sbuf_p0_rdat_1039 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1040 = {_zz_shareBuffer_sbuf_p0_rdat_1041,_zz_shareBuffer_sbuf_p0_rdat_1042};
  assign _zz_shareBuffer_sbuf_p0_rdat_1153 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1154 = {_zz_shareBuffer_sbuf_p0_rdat_1155,_zz_shareBuffer_sbuf_p0_rdat_1156};
  assign _zz_shareBuffer_sbuf_p0_rdat_1266 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1267 = {_zz_shareBuffer_sbuf_p0_rdat_1268,_zz_shareBuffer_sbuf_p0_rdat_1269};
  assign _zz_shareBuffer_sbuf_p0_rdat_1379 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1380 = {_zz_shareBuffer_sbuf_p0_rdat_1381,_zz_shareBuffer_sbuf_p0_rdat_1382};
  assign _zz_shareBuffer_sbuf_p0_rdat_1491 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1492 = {_zz_shareBuffer_sbuf_p0_rdat_1493,_zz_shareBuffer_sbuf_p0_rdat_1494};
  assign _zz_shareBuffer_sbuf_p0_rdat_1603 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1604 = {_zz_shareBuffer_sbuf_p0_rdat_1605,_zz_shareBuffer_sbuf_p0_rdat_1606};
  assign _zz_shareBuffer_sbuf_p0_rdat_1713 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1714 = {_zz_shareBuffer_sbuf_p0_rdat_1715,_zz_shareBuffer_sbuf_p0_rdat_1716};
  assign _zz_shareBuffer_sbuf_p0_rdat_30 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_31 = {_zz_shareBuffer_sbuf_p0_rdat_32,_zz_shareBuffer_sbuf_p0_rdat_33};
  assign _zz_shareBuffer_sbuf_p0_rdat_139 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_140 = {_zz_shareBuffer_sbuf_p0_rdat_141,_zz_shareBuffer_sbuf_p0_rdat_142};
  assign _zz_shareBuffer_sbuf_p0_rdat_250 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_251 = {_zz_shareBuffer_sbuf_p0_rdat_252,_zz_shareBuffer_sbuf_p0_rdat_253};
  assign _zz_shareBuffer_sbuf_p0_rdat_361 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_362 = {_zz_shareBuffer_sbuf_p0_rdat_363,_zz_shareBuffer_sbuf_p0_rdat_364};
  assign _zz_shareBuffer_sbuf_p0_rdat_474 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_475 = {_zz_shareBuffer_sbuf_p0_rdat_476,_zz_shareBuffer_sbuf_p0_rdat_477};
  assign _zz_shareBuffer_sbuf_p0_rdat_587 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_588 = {_zz_shareBuffer_sbuf_p0_rdat_589,_zz_shareBuffer_sbuf_p0_rdat_590};
  assign _zz_shareBuffer_sbuf_p0_rdat_700 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_701 = {_zz_shareBuffer_sbuf_p0_rdat_702,_zz_shareBuffer_sbuf_p0_rdat_703};
  assign _zz_shareBuffer_sbuf_p0_rdat_813 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_814 = {_zz_shareBuffer_sbuf_p0_rdat_815,_zz_shareBuffer_sbuf_p0_rdat_816};
  assign _zz_shareBuffer_sbuf_p0_rdat_928 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_929 = {_zz_shareBuffer_sbuf_p0_rdat_930,_zz_shareBuffer_sbuf_p0_rdat_931};
  assign _zz_shareBuffer_sbuf_p0_rdat_1041 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1042 = {_zz_shareBuffer_sbuf_p0_rdat_1043,_zz_shareBuffer_sbuf_p0_rdat_1044};
  assign _zz_shareBuffer_sbuf_p0_rdat_1155 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1156 = {_zz_shareBuffer_sbuf_p0_rdat_1157,_zz_shareBuffer_sbuf_p0_rdat_1158};
  assign _zz_shareBuffer_sbuf_p0_rdat_1268 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1269 = {_zz_shareBuffer_sbuf_p0_rdat_1270,_zz_shareBuffer_sbuf_p0_rdat_1271};
  assign _zz_shareBuffer_sbuf_p0_rdat_1381 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1382 = {_zz_shareBuffer_sbuf_p0_rdat_1383,_zz_shareBuffer_sbuf_p0_rdat_1384};
  assign _zz_shareBuffer_sbuf_p0_rdat_1493 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1494 = {_zz_shareBuffer_sbuf_p0_rdat_1495,_zz_shareBuffer_sbuf_p0_rdat_1496};
  assign _zz_shareBuffer_sbuf_p0_rdat_1605 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1606 = {_zz_shareBuffer_sbuf_p0_rdat_1607,_zz_shareBuffer_sbuf_p0_rdat_1608};
  assign _zz_shareBuffer_sbuf_p0_rdat_1715 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1716 = {_zz_shareBuffer_sbuf_p0_rdat_1717,_zz_shareBuffer_sbuf_p0_rdat_1718};
  assign _zz_shareBuffer_sbuf_p0_rdat_32 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_33 = {_zz_shareBuffer_sbuf_p0_rdat_34,_zz_shareBuffer_sbuf_p0_rdat_35};
  assign _zz_shareBuffer_sbuf_p0_rdat_141 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_142 = {_zz_shareBuffer_sbuf_p0_rdat_143,_zz_shareBuffer_sbuf_p0_rdat_144};
  assign _zz_shareBuffer_sbuf_p0_rdat_252 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_253 = {_zz_shareBuffer_sbuf_p0_rdat_254,_zz_shareBuffer_sbuf_p0_rdat_255};
  assign _zz_shareBuffer_sbuf_p0_rdat_363 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_364 = {_zz_shareBuffer_sbuf_p0_rdat_365,_zz_shareBuffer_sbuf_p0_rdat_366};
  assign _zz_shareBuffer_sbuf_p0_rdat_476 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_477 = {_zz_shareBuffer_sbuf_p0_rdat_478,_zz_shareBuffer_sbuf_p0_rdat_479};
  assign _zz_shareBuffer_sbuf_p0_rdat_589 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_590 = {_zz_shareBuffer_sbuf_p0_rdat_591,_zz_shareBuffer_sbuf_p0_rdat_592};
  assign _zz_shareBuffer_sbuf_p0_rdat_702 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_703 = {_zz_shareBuffer_sbuf_p0_rdat_704,_zz_shareBuffer_sbuf_p0_rdat_705};
  assign _zz_shareBuffer_sbuf_p0_rdat_815 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_816 = {_zz_shareBuffer_sbuf_p0_rdat_817,_zz_shareBuffer_sbuf_p0_rdat_818};
  assign _zz_shareBuffer_sbuf_p0_rdat_930 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_931 = {_zz_shareBuffer_sbuf_p0_rdat_932,_zz_shareBuffer_sbuf_p0_rdat_933};
  assign _zz_shareBuffer_sbuf_p0_rdat_1043 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1044 = {_zz_shareBuffer_sbuf_p0_rdat_1045,_zz_shareBuffer_sbuf_p0_rdat_1046};
  assign _zz_shareBuffer_sbuf_p0_rdat_1157 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1158 = {_zz_shareBuffer_sbuf_p0_rdat_1159,_zz_shareBuffer_sbuf_p0_rdat_1160};
  assign _zz_shareBuffer_sbuf_p0_rdat_1270 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1271 = {_zz_shareBuffer_sbuf_p0_rdat_1272,_zz_shareBuffer_sbuf_p0_rdat_1273};
  assign _zz_shareBuffer_sbuf_p0_rdat_1383 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1384 = {_zz_shareBuffer_sbuf_p0_rdat_1385,_zz_shareBuffer_sbuf_p0_rdat_1386};
  assign _zz_shareBuffer_sbuf_p0_rdat_1495 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1496 = {_zz_shareBuffer_sbuf_p0_rdat_1497,_zz_shareBuffer_sbuf_p0_rdat_1498};
  assign _zz_shareBuffer_sbuf_p0_rdat_1607 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1608 = {_zz_shareBuffer_sbuf_p0_rdat_1609,_zz_shareBuffer_sbuf_p0_rdat_1610};
  assign _zz_shareBuffer_sbuf_p0_rdat_1717 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1718 = {_zz_shareBuffer_sbuf_p0_rdat_1719,_zz_shareBuffer_sbuf_p0_rdat_1720};
  assign _zz_shareBuffer_sbuf_p0_rdat_34 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_35 = {_zz_shareBuffer_sbuf_p0_rdat_36,_zz_shareBuffer_sbuf_p0_rdat_37};
  assign _zz_shareBuffer_sbuf_p0_rdat_143 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_144 = {_zz_shareBuffer_sbuf_p0_rdat_145,_zz_shareBuffer_sbuf_p0_rdat_146};
  assign _zz_shareBuffer_sbuf_p0_rdat_254 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_255 = {_zz_shareBuffer_sbuf_p0_rdat_256,_zz_shareBuffer_sbuf_p0_rdat_257};
  assign _zz_shareBuffer_sbuf_p0_rdat_365 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_366 = {_zz_shareBuffer_sbuf_p0_rdat_367,_zz_shareBuffer_sbuf_p0_rdat_368};
  assign _zz_shareBuffer_sbuf_p0_rdat_478 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_479 = {_zz_shareBuffer_sbuf_p0_rdat_480,_zz_shareBuffer_sbuf_p0_rdat_481};
  assign _zz_shareBuffer_sbuf_p0_rdat_591 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_592 = {_zz_shareBuffer_sbuf_p0_rdat_593,_zz_shareBuffer_sbuf_p0_rdat_594};
  assign _zz_shareBuffer_sbuf_p0_rdat_704 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_705 = {_zz_shareBuffer_sbuf_p0_rdat_706,_zz_shareBuffer_sbuf_p0_rdat_707};
  assign _zz_shareBuffer_sbuf_p0_rdat_817 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_818 = {_zz_shareBuffer_sbuf_p0_rdat_819,_zz_shareBuffer_sbuf_p0_rdat_820};
  assign _zz_shareBuffer_sbuf_p0_rdat_932 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_933 = {_zz_shareBuffer_sbuf_p0_rdat_934,_zz_shareBuffer_sbuf_p0_rdat_935};
  assign _zz_shareBuffer_sbuf_p0_rdat_1045 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1046 = {_zz_shareBuffer_sbuf_p0_rdat_1047,_zz_shareBuffer_sbuf_p0_rdat_1048};
  assign _zz_shareBuffer_sbuf_p0_rdat_1159 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1160 = {_zz_shareBuffer_sbuf_p0_rdat_1161,_zz_shareBuffer_sbuf_p0_rdat_1162};
  assign _zz_shareBuffer_sbuf_p0_rdat_1272 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1273 = {_zz_shareBuffer_sbuf_p0_rdat_1274,_zz_shareBuffer_sbuf_p0_rdat_1275};
  assign _zz_shareBuffer_sbuf_p0_rdat_1385 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1386 = {_zz_shareBuffer_sbuf_p0_rdat_1387,_zz_shareBuffer_sbuf_p0_rdat_1388};
  assign _zz_shareBuffer_sbuf_p0_rdat_1497 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1498 = {_zz_shareBuffer_sbuf_p0_rdat_1499,_zz_shareBuffer_sbuf_p0_rdat_1500};
  assign _zz_shareBuffer_sbuf_p0_rdat_1609 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1610 = {_zz_shareBuffer_sbuf_p0_rdat_1611,_zz_shareBuffer_sbuf_p0_rdat_1612};
  assign _zz_shareBuffer_sbuf_p0_rdat_1719 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1720 = {_zz_shareBuffer_sbuf_p0_rdat_1721,_zz_shareBuffer_sbuf_p0_rdat_1722};
  assign _zz_shareBuffer_sbuf_p0_rdat_36 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_37 = {_zz_shareBuffer_sbuf_p0_rdat_38,_zz_shareBuffer_sbuf_p0_rdat_39};
  assign _zz_shareBuffer_sbuf_p0_rdat_145 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_146 = {_zz_shareBuffer_sbuf_p0_rdat_147,_zz_shareBuffer_sbuf_p0_rdat_148};
  assign _zz_shareBuffer_sbuf_p0_rdat_256 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_257 = {_zz_shareBuffer_sbuf_p0_rdat_258,_zz_shareBuffer_sbuf_p0_rdat_259};
  assign _zz_shareBuffer_sbuf_p0_rdat_367 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_368 = {_zz_shareBuffer_sbuf_p0_rdat_369,_zz_shareBuffer_sbuf_p0_rdat_370};
  assign _zz_shareBuffer_sbuf_p0_rdat_480 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_481 = {_zz_shareBuffer_sbuf_p0_rdat_482,_zz_shareBuffer_sbuf_p0_rdat_483};
  assign _zz_shareBuffer_sbuf_p0_rdat_593 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_594 = {_zz_shareBuffer_sbuf_p0_rdat_595,_zz_shareBuffer_sbuf_p0_rdat_596};
  assign _zz_shareBuffer_sbuf_p0_rdat_706 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_707 = {_zz_shareBuffer_sbuf_p0_rdat_708,_zz_shareBuffer_sbuf_p0_rdat_709};
  assign _zz_shareBuffer_sbuf_p0_rdat_819 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_820 = {_zz_shareBuffer_sbuf_p0_rdat_821,_zz_shareBuffer_sbuf_p0_rdat_822};
  assign _zz_shareBuffer_sbuf_p0_rdat_934 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_935 = {_zz_shareBuffer_sbuf_p0_rdat_936,_zz_shareBuffer_sbuf_p0_rdat_937};
  assign _zz_shareBuffer_sbuf_p0_rdat_1047 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1048 = {_zz_shareBuffer_sbuf_p0_rdat_1049,_zz_shareBuffer_sbuf_p0_rdat_1050};
  assign _zz_shareBuffer_sbuf_p0_rdat_1161 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1162 = {_zz_shareBuffer_sbuf_p0_rdat_1163,_zz_shareBuffer_sbuf_p0_rdat_1164};
  assign _zz_shareBuffer_sbuf_p0_rdat_1274 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1275 = {_zz_shareBuffer_sbuf_p0_rdat_1276,_zz_shareBuffer_sbuf_p0_rdat_1277};
  assign _zz_shareBuffer_sbuf_p0_rdat_1387 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1388 = {_zz_shareBuffer_sbuf_p0_rdat_1389,_zz_shareBuffer_sbuf_p0_rdat_1390};
  assign _zz_shareBuffer_sbuf_p0_rdat_1499 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1500 = {_zz_shareBuffer_sbuf_p0_rdat_1501,_zz_shareBuffer_sbuf_p0_rdat_1502};
  assign _zz_shareBuffer_sbuf_p0_rdat_1611 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1612 = {_zz_shareBuffer_sbuf_p0_rdat_1613,_zz_shareBuffer_sbuf_p0_rdat_1614};
  assign _zz_shareBuffer_sbuf_p0_rdat_1721 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1722 = {_zz_shareBuffer_sbuf_p0_rdat_1723,_zz_shareBuffer_sbuf_p0_rdat_1724};
  assign _zz_shareBuffer_sbuf_p0_rdat_38 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_39 = {_zz_shareBuffer_sbuf_p0_rdat_40,_zz_shareBuffer_sbuf_p0_rdat_41};
  assign _zz_shareBuffer_sbuf_p0_rdat_147 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_148 = {_zz_shareBuffer_sbuf_p0_rdat_149,_zz_shareBuffer_sbuf_p0_rdat_150};
  assign _zz_shareBuffer_sbuf_p0_rdat_258 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_259 = {_zz_shareBuffer_sbuf_p0_rdat_260,_zz_shareBuffer_sbuf_p0_rdat_261};
  assign _zz_shareBuffer_sbuf_p0_rdat_369 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_370 = {_zz_shareBuffer_sbuf_p0_rdat_371,_zz_shareBuffer_sbuf_p0_rdat_372};
  assign _zz_shareBuffer_sbuf_p0_rdat_482 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_483 = {_zz_shareBuffer_sbuf_p0_rdat_484,_zz_shareBuffer_sbuf_p0_rdat_485};
  assign _zz_shareBuffer_sbuf_p0_rdat_595 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_596 = {_zz_shareBuffer_sbuf_p0_rdat_597,_zz_shareBuffer_sbuf_p0_rdat_598};
  assign _zz_shareBuffer_sbuf_p0_rdat_708 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_709 = {_zz_shareBuffer_sbuf_p0_rdat_710,_zz_shareBuffer_sbuf_p0_rdat_711};
  assign _zz_shareBuffer_sbuf_p0_rdat_821 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_822 = {_zz_shareBuffer_sbuf_p0_rdat_823,_zz_shareBuffer_sbuf_p0_rdat_824};
  assign _zz_shareBuffer_sbuf_p0_rdat_936 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_937 = {_zz_shareBuffer_sbuf_p0_rdat_938,_zz_shareBuffer_sbuf_p0_rdat_939};
  assign _zz_shareBuffer_sbuf_p0_rdat_1049 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1050 = {_zz_shareBuffer_sbuf_p0_rdat_1051,_zz_shareBuffer_sbuf_p0_rdat_1052};
  assign _zz_shareBuffer_sbuf_p0_rdat_1163 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1164 = {_zz_shareBuffer_sbuf_p0_rdat_1165,_zz_shareBuffer_sbuf_p0_rdat_1166};
  assign _zz_shareBuffer_sbuf_p0_rdat_1276 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1277 = {_zz_shareBuffer_sbuf_p0_rdat_1278,_zz_shareBuffer_sbuf_p0_rdat_1279};
  assign _zz_shareBuffer_sbuf_p0_rdat_1389 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1390 = {_zz_shareBuffer_sbuf_p0_rdat_1391,_zz_shareBuffer_sbuf_p0_rdat_1392};
  assign _zz_shareBuffer_sbuf_p0_rdat_1501 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1502 = {_zz_shareBuffer_sbuf_p0_rdat_1503,_zz_shareBuffer_sbuf_p0_rdat_1504};
  assign _zz_shareBuffer_sbuf_p0_rdat_1613 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1614 = {_zz_shareBuffer_sbuf_p0_rdat_1615,_zz_shareBuffer_sbuf_p0_rdat_1616};
  assign _zz_shareBuffer_sbuf_p0_rdat_1723 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1724 = {_zz_shareBuffer_sbuf_p0_rdat_1725,_zz_shareBuffer_sbuf_p0_rdat_1726};
  assign _zz_shareBuffer_sbuf_p0_rdat_40 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_41 = {_zz_shareBuffer_sbuf_p0_rdat_42,_zz_shareBuffer_sbuf_p0_rdat_43};
  assign _zz_shareBuffer_sbuf_p0_rdat_149 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_150 = {_zz_shareBuffer_sbuf_p0_rdat_151,_zz_shareBuffer_sbuf_p0_rdat_152};
  assign _zz_shareBuffer_sbuf_p0_rdat_260 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_261 = {_zz_shareBuffer_sbuf_p0_rdat_262,_zz_shareBuffer_sbuf_p0_rdat_263};
  assign _zz_shareBuffer_sbuf_p0_rdat_371 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_372 = {_zz_shareBuffer_sbuf_p0_rdat_373,_zz_shareBuffer_sbuf_p0_rdat_374};
  assign _zz_shareBuffer_sbuf_p0_rdat_484 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_485 = {_zz_shareBuffer_sbuf_p0_rdat_486,_zz_shareBuffer_sbuf_p0_rdat_487};
  assign _zz_shareBuffer_sbuf_p0_rdat_597 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_598 = {_zz_shareBuffer_sbuf_p0_rdat_599,_zz_shareBuffer_sbuf_p0_rdat_600};
  assign _zz_shareBuffer_sbuf_p0_rdat_710 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_711 = {_zz_shareBuffer_sbuf_p0_rdat_712,_zz_shareBuffer_sbuf_p0_rdat_713};
  assign _zz_shareBuffer_sbuf_p0_rdat_823 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_824 = {_zz_shareBuffer_sbuf_p0_rdat_825,_zz_shareBuffer_sbuf_p0_rdat_826};
  assign _zz_shareBuffer_sbuf_p0_rdat_938 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_939 = {_zz_shareBuffer_sbuf_p0_rdat_940,_zz_shareBuffer_sbuf_p0_rdat_941};
  assign _zz_shareBuffer_sbuf_p0_rdat_1051 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1052 = {_zz_shareBuffer_sbuf_p0_rdat_1053,_zz_shareBuffer_sbuf_p0_rdat_1054};
  assign _zz_shareBuffer_sbuf_p0_rdat_1165 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1166 = {_zz_shareBuffer_sbuf_p0_rdat_1167,_zz_shareBuffer_sbuf_p0_rdat_1168};
  assign _zz_shareBuffer_sbuf_p0_rdat_1278 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1279 = {_zz_shareBuffer_sbuf_p0_rdat_1280,_zz_shareBuffer_sbuf_p0_rdat_1281};
  assign _zz_shareBuffer_sbuf_p0_rdat_1391 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1392 = {_zz_shareBuffer_sbuf_p0_rdat_1393,_zz_shareBuffer_sbuf_p0_rdat_1394};
  assign _zz_shareBuffer_sbuf_p0_rdat_1503 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1504 = {_zz_shareBuffer_sbuf_p0_rdat_1505,_zz_shareBuffer_sbuf_p0_rdat_1506};
  assign _zz_shareBuffer_sbuf_p0_rdat_1615 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1616 = {_zz_shareBuffer_sbuf_p0_rdat_1617,_zz_shareBuffer_sbuf_p0_rdat_1618};
  assign _zz_shareBuffer_sbuf_p0_rdat_1725 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1726 = {_zz_shareBuffer_sbuf_p0_rdat_1727,_zz_shareBuffer_sbuf_p0_rdat_1728};
  assign _zz_shareBuffer_sbuf_p0_rdat_42 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_43 = {_zz_shareBuffer_sbuf_p0_rdat_44,_zz_shareBuffer_sbuf_p0_rdat_45};
  assign _zz_shareBuffer_sbuf_p0_rdat_151 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_152 = {_zz_shareBuffer_sbuf_p0_rdat_153,_zz_shareBuffer_sbuf_p0_rdat_154};
  assign _zz_shareBuffer_sbuf_p0_rdat_262 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_263 = {_zz_shareBuffer_sbuf_p0_rdat_264,_zz_shareBuffer_sbuf_p0_rdat_265};
  assign _zz_shareBuffer_sbuf_p0_rdat_373 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_374 = {_zz_shareBuffer_sbuf_p0_rdat_375,_zz_shareBuffer_sbuf_p0_rdat_376};
  assign _zz_shareBuffer_sbuf_p0_rdat_486 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_487 = {_zz_shareBuffer_sbuf_p0_rdat_488,_zz_shareBuffer_sbuf_p0_rdat_489};
  assign _zz_shareBuffer_sbuf_p0_rdat_599 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_600 = {_zz_shareBuffer_sbuf_p0_rdat_601,_zz_shareBuffer_sbuf_p0_rdat_602};
  assign _zz_shareBuffer_sbuf_p0_rdat_712 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_713 = {_zz_shareBuffer_sbuf_p0_rdat_714,_zz_shareBuffer_sbuf_p0_rdat_715};
  assign _zz_shareBuffer_sbuf_p0_rdat_825 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_826 = {_zz_shareBuffer_sbuf_p0_rdat_827,_zz_shareBuffer_sbuf_p0_rdat_828};
  assign _zz_shareBuffer_sbuf_p0_rdat_940 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_941 = {_zz_shareBuffer_sbuf_p0_rdat_942,_zz_shareBuffer_sbuf_p0_rdat_943};
  assign _zz_shareBuffer_sbuf_p0_rdat_1053 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1054 = {_zz_shareBuffer_sbuf_p0_rdat_1055,_zz_shareBuffer_sbuf_p0_rdat_1056};
  assign _zz_shareBuffer_sbuf_p0_rdat_1167 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1168 = {_zz_shareBuffer_sbuf_p0_rdat_1169,_zz_shareBuffer_sbuf_p0_rdat_1170};
  assign _zz_shareBuffer_sbuf_p0_rdat_1280 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1281 = {_zz_shareBuffer_sbuf_p0_rdat_1282,_zz_shareBuffer_sbuf_p0_rdat_1283};
  assign _zz_shareBuffer_sbuf_p0_rdat_1393 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1394 = {_zz_shareBuffer_sbuf_p0_rdat_1395,_zz_shareBuffer_sbuf_p0_rdat_1396};
  assign _zz_shareBuffer_sbuf_p0_rdat_1505 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1506 = {_zz_shareBuffer_sbuf_p0_rdat_1507,_zz_shareBuffer_sbuf_p0_rdat_1508};
  assign _zz_shareBuffer_sbuf_p0_rdat_1617 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1618 = {_zz_shareBuffer_sbuf_p0_rdat_1619,_zz_shareBuffer_sbuf_p0_rdat_1620};
  assign _zz_shareBuffer_sbuf_p0_rdat_1727 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1728 = {_zz_shareBuffer_sbuf_p0_rdat_1729,_zz_shareBuffer_sbuf_p0_rdat_1730};
  assign _zz_shareBuffer_sbuf_p0_rdat_44 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_45 = {_zz_shareBuffer_sbuf_p0_rdat_46,_zz_shareBuffer_sbuf_p0_rdat_47};
  assign _zz_shareBuffer_sbuf_p0_rdat_153 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_154 = {_zz_shareBuffer_sbuf_p0_rdat_155,_zz_shareBuffer_sbuf_p0_rdat_156};
  assign _zz_shareBuffer_sbuf_p0_rdat_264 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_265 = {_zz_shareBuffer_sbuf_p0_rdat_266,_zz_shareBuffer_sbuf_p0_rdat_267};
  assign _zz_shareBuffer_sbuf_p0_rdat_375 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_376 = {_zz_shareBuffer_sbuf_p0_rdat_377,_zz_shareBuffer_sbuf_p0_rdat_378};
  assign _zz_shareBuffer_sbuf_p0_rdat_488 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_489 = {_zz_shareBuffer_sbuf_p0_rdat_490,_zz_shareBuffer_sbuf_p0_rdat_491};
  assign _zz_shareBuffer_sbuf_p0_rdat_601 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_602 = {_zz_shareBuffer_sbuf_p0_rdat_603,_zz_shareBuffer_sbuf_p0_rdat_604};
  assign _zz_shareBuffer_sbuf_p0_rdat_714 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_715 = {_zz_shareBuffer_sbuf_p0_rdat_716,_zz_shareBuffer_sbuf_p0_rdat_717};
  assign _zz_shareBuffer_sbuf_p0_rdat_827 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_828 = {_zz_shareBuffer_sbuf_p0_rdat_829,_zz_shareBuffer_sbuf_p0_rdat_830};
  assign _zz_shareBuffer_sbuf_p0_rdat_942 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_943 = {_zz_shareBuffer_sbuf_p0_rdat_944,_zz_shareBuffer_sbuf_p0_rdat_945};
  assign _zz_shareBuffer_sbuf_p0_rdat_1055 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1056 = {_zz_shareBuffer_sbuf_p0_rdat_1057,_zz_shareBuffer_sbuf_p0_rdat_1058};
  assign _zz_shareBuffer_sbuf_p0_rdat_1169 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1170 = {_zz_shareBuffer_sbuf_p0_rdat_1171,_zz_shareBuffer_sbuf_p0_rdat_1172};
  assign _zz_shareBuffer_sbuf_p0_rdat_1282 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1283 = {_zz_shareBuffer_sbuf_p0_rdat_1284,_zz_shareBuffer_sbuf_p0_rdat_1285};
  assign _zz_shareBuffer_sbuf_p0_rdat_1395 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1396 = {_zz_shareBuffer_sbuf_p0_rdat_1397,_zz_shareBuffer_sbuf_p0_rdat_1398};
  assign _zz_shareBuffer_sbuf_p0_rdat_1507 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1508 = {_zz_shareBuffer_sbuf_p0_rdat_1509,_zz_shareBuffer_sbuf_p0_rdat_1510};
  assign _zz_shareBuffer_sbuf_p0_rdat_1619 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1620 = {_zz_shareBuffer_sbuf_p0_rdat_1621,_zz_shareBuffer_sbuf_p0_rdat_1622};
  assign _zz_shareBuffer_sbuf_p0_rdat_1729 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1730 = {_zz_shareBuffer_sbuf_p0_rdat_1731,_zz_shareBuffer_sbuf_p0_rdat_1732};
  assign _zz_shareBuffer_sbuf_p0_rdat_46 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_47 = {_zz_shareBuffer_sbuf_p0_rdat_48,_zz_shareBuffer_sbuf_p0_rdat_49};
  assign _zz_shareBuffer_sbuf_p0_rdat_155 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_156 = {_zz_shareBuffer_sbuf_p0_rdat_157,_zz_shareBuffer_sbuf_p0_rdat_158};
  assign _zz_shareBuffer_sbuf_p0_rdat_266 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_267 = {_zz_shareBuffer_sbuf_p0_rdat_268,_zz_shareBuffer_sbuf_p0_rdat_269};
  assign _zz_shareBuffer_sbuf_p0_rdat_377 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_378 = {_zz_shareBuffer_sbuf_p0_rdat_379,_zz_shareBuffer_sbuf_p0_rdat_380};
  assign _zz_shareBuffer_sbuf_p0_rdat_490 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_491 = {_zz_shareBuffer_sbuf_p0_rdat_492,_zz_shareBuffer_sbuf_p0_rdat_493};
  assign _zz_shareBuffer_sbuf_p0_rdat_603 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_604 = {_zz_shareBuffer_sbuf_p0_rdat_605,_zz_shareBuffer_sbuf_p0_rdat_606};
  assign _zz_shareBuffer_sbuf_p0_rdat_716 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_717 = {_zz_shareBuffer_sbuf_p0_rdat_718,_zz_shareBuffer_sbuf_p0_rdat_719};
  assign _zz_shareBuffer_sbuf_p0_rdat_829 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_830 = {_zz_shareBuffer_sbuf_p0_rdat_831,_zz_shareBuffer_sbuf_p0_rdat_832};
  assign _zz_shareBuffer_sbuf_p0_rdat_944 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_945 = {_zz_shareBuffer_sbuf_p0_rdat_946,_zz_shareBuffer_sbuf_p0_rdat_947};
  assign _zz_shareBuffer_sbuf_p0_rdat_1057 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1058 = {_zz_shareBuffer_sbuf_p0_rdat_1059,_zz_shareBuffer_sbuf_p0_rdat_1060};
  assign _zz_shareBuffer_sbuf_p0_rdat_1171 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1172 = {_zz_shareBuffer_sbuf_p0_rdat_1173,_zz_shareBuffer_sbuf_p0_rdat_1174};
  assign _zz_shareBuffer_sbuf_p0_rdat_1284 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1285 = {_zz_shareBuffer_sbuf_p0_rdat_1286,_zz_shareBuffer_sbuf_p0_rdat_1287};
  assign _zz_shareBuffer_sbuf_p0_rdat_1397 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1398 = {_zz_shareBuffer_sbuf_p0_rdat_1399,_zz_shareBuffer_sbuf_p0_rdat_1400};
  assign _zz_shareBuffer_sbuf_p0_rdat_1509 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1510 = {_zz_shareBuffer_sbuf_p0_rdat_1511,_zz_shareBuffer_sbuf_p0_rdat_1512};
  assign _zz_shareBuffer_sbuf_p0_rdat_1621 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1622 = {_zz_shareBuffer_sbuf_p0_rdat_1623,_zz_shareBuffer_sbuf_p0_rdat_1624};
  assign _zz_shareBuffer_sbuf_p0_rdat_1731 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1732 = {_zz_shareBuffer_sbuf_p0_rdat_1733,_zz_shareBuffer_sbuf_p0_rdat_1734};
  assign _zz_shareBuffer_sbuf_p0_rdat_48 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_49 = {_zz_shareBuffer_sbuf_p0_rdat_50,_zz_shareBuffer_sbuf_p0_rdat_51};
  assign _zz_shareBuffer_sbuf_p0_rdat_157 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_158 = {_zz_shareBuffer_sbuf_p0_rdat_159,_zz_shareBuffer_sbuf_p0_rdat_160};
  assign _zz_shareBuffer_sbuf_p0_rdat_268 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_269 = {_zz_shareBuffer_sbuf_p0_rdat_270,_zz_shareBuffer_sbuf_p0_rdat_271};
  assign _zz_shareBuffer_sbuf_p0_rdat_379 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_380 = {_zz_shareBuffer_sbuf_p0_rdat_381,_zz_shareBuffer_sbuf_p0_rdat_382};
  assign _zz_shareBuffer_sbuf_p0_rdat_492 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_493 = {_zz_shareBuffer_sbuf_p0_rdat_494,_zz_shareBuffer_sbuf_p0_rdat_495};
  assign _zz_shareBuffer_sbuf_p0_rdat_605 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_606 = {_zz_shareBuffer_sbuf_p0_rdat_607,_zz_shareBuffer_sbuf_p0_rdat_608};
  assign _zz_shareBuffer_sbuf_p0_rdat_718 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_719 = {_zz_shareBuffer_sbuf_p0_rdat_720,_zz_shareBuffer_sbuf_p0_rdat_721};
  assign _zz_shareBuffer_sbuf_p0_rdat_831 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_832 = {_zz_shareBuffer_sbuf_p0_rdat_833,_zz_shareBuffer_sbuf_p0_rdat_834};
  assign _zz_shareBuffer_sbuf_p0_rdat_946 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_947 = {_zz_shareBuffer_sbuf_p0_rdat_948,_zz_shareBuffer_sbuf_p0_rdat_949};
  assign _zz_shareBuffer_sbuf_p0_rdat_1059 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1060 = {_zz_shareBuffer_sbuf_p0_rdat_1061,_zz_shareBuffer_sbuf_p0_rdat_1062};
  assign _zz_shareBuffer_sbuf_p0_rdat_1173 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1174 = {_zz_shareBuffer_sbuf_p0_rdat_1175,_zz_shareBuffer_sbuf_p0_rdat_1176};
  assign _zz_shareBuffer_sbuf_p0_rdat_1286 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1287 = {_zz_shareBuffer_sbuf_p0_rdat_1288,_zz_shareBuffer_sbuf_p0_rdat_1289};
  assign _zz_shareBuffer_sbuf_p0_rdat_1399 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1400 = {_zz_shareBuffer_sbuf_p0_rdat_1401,_zz_shareBuffer_sbuf_p0_rdat_1402};
  assign _zz_shareBuffer_sbuf_p0_rdat_1511 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1512 = {_zz_shareBuffer_sbuf_p0_rdat_1513,_zz_shareBuffer_sbuf_p0_rdat_1514};
  assign _zz_shareBuffer_sbuf_p0_rdat_1623 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1624 = {_zz_shareBuffer_sbuf_p0_rdat_1625,_zz_shareBuffer_sbuf_p0_rdat_1626};
  assign _zz_shareBuffer_sbuf_p0_rdat_1733 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1734 = {_zz_shareBuffer_sbuf_p0_rdat_1735,_zz_shareBuffer_sbuf_p0_rdat_1736};
  assign _zz_shareBuffer_sbuf_p0_rdat_50 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_51 = {_zz_shareBuffer_sbuf_p0_rdat_52,_zz_shareBuffer_sbuf_p0_rdat_53};
  assign _zz_shareBuffer_sbuf_p0_rdat_159 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_160 = {_zz_shareBuffer_sbuf_p0_rdat_161,_zz_shareBuffer_sbuf_p0_rdat_162};
  assign _zz_shareBuffer_sbuf_p0_rdat_270 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_271 = {_zz_shareBuffer_sbuf_p0_rdat_272,_zz_shareBuffer_sbuf_p0_rdat_273};
  assign _zz_shareBuffer_sbuf_p0_rdat_381 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_382 = {_zz_shareBuffer_sbuf_p0_rdat_383,_zz_shareBuffer_sbuf_p0_rdat_384};
  assign _zz_shareBuffer_sbuf_p0_rdat_494 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_495 = {_zz_shareBuffer_sbuf_p0_rdat_496,_zz_shareBuffer_sbuf_p0_rdat_497};
  assign _zz_shareBuffer_sbuf_p0_rdat_607 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_608 = {_zz_shareBuffer_sbuf_p0_rdat_609,_zz_shareBuffer_sbuf_p0_rdat_610};
  assign _zz_shareBuffer_sbuf_p0_rdat_720 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_721 = {_zz_shareBuffer_sbuf_p0_rdat_722,_zz_shareBuffer_sbuf_p0_rdat_723};
  assign _zz_shareBuffer_sbuf_p0_rdat_833 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_834 = {_zz_shareBuffer_sbuf_p0_rdat_835,_zz_shareBuffer_sbuf_p0_rdat_836};
  assign _zz_shareBuffer_sbuf_p0_rdat_948 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_949 = {_zz_shareBuffer_sbuf_p0_rdat_950,_zz_shareBuffer_sbuf_p0_rdat_951};
  assign _zz_shareBuffer_sbuf_p0_rdat_1061 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1062 = {_zz_shareBuffer_sbuf_p0_rdat_1063,_zz_shareBuffer_sbuf_p0_rdat_1064};
  assign _zz_shareBuffer_sbuf_p0_rdat_1175 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1176 = {_zz_shareBuffer_sbuf_p0_rdat_1177,_zz_shareBuffer_sbuf_p0_rdat_1178};
  assign _zz_shareBuffer_sbuf_p0_rdat_1288 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1289 = {_zz_shareBuffer_sbuf_p0_rdat_1290,_zz_shareBuffer_sbuf_p0_rdat_1291};
  assign _zz_shareBuffer_sbuf_p0_rdat_1401 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1402 = {_zz_shareBuffer_sbuf_p0_rdat_1403,_zz_shareBuffer_sbuf_p0_rdat_1404};
  assign _zz_shareBuffer_sbuf_p0_rdat_1513 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1514 = {_zz_shareBuffer_sbuf_p0_rdat_1515,_zz_shareBuffer_sbuf_p0_rdat_1516};
  assign _zz_shareBuffer_sbuf_p0_rdat_1625 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1626 = {_zz_shareBuffer_sbuf_p0_rdat_1627,_zz_shareBuffer_sbuf_p0_rdat_1628};
  assign _zz_shareBuffer_sbuf_p0_rdat_1735 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1736 = {_zz_shareBuffer_sbuf_p0_rdat_1737,_zz_shareBuffer_sbuf_p0_rdat_1738};
  assign _zz_shareBuffer_sbuf_p0_rdat_52 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_53 = {_zz_shareBuffer_sbuf_p0_rdat_54,_zz_shareBuffer_sbuf_p0_rdat_55};
  assign _zz_shareBuffer_sbuf_p0_rdat_161 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_162 = {_zz_shareBuffer_sbuf_p0_rdat_163,_zz_shareBuffer_sbuf_p0_rdat_164};
  assign _zz_shareBuffer_sbuf_p0_rdat_272 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_273 = {_zz_shareBuffer_sbuf_p0_rdat_274,_zz_shareBuffer_sbuf_p0_rdat_275};
  assign _zz_shareBuffer_sbuf_p0_rdat_383 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_384 = {_zz_shareBuffer_sbuf_p0_rdat_385,_zz_shareBuffer_sbuf_p0_rdat_386};
  assign _zz_shareBuffer_sbuf_p0_rdat_496 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_497 = {_zz_shareBuffer_sbuf_p0_rdat_498,_zz_shareBuffer_sbuf_p0_rdat_499};
  assign _zz_shareBuffer_sbuf_p0_rdat_609 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_610 = {_zz_shareBuffer_sbuf_p0_rdat_611,_zz_shareBuffer_sbuf_p0_rdat_612};
  assign _zz_shareBuffer_sbuf_p0_rdat_722 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_723 = {_zz_shareBuffer_sbuf_p0_rdat_724,_zz_shareBuffer_sbuf_p0_rdat_725};
  assign _zz_shareBuffer_sbuf_p0_rdat_835 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_836 = {_zz_shareBuffer_sbuf_p0_rdat_837,_zz_shareBuffer_sbuf_p0_rdat_838};
  assign _zz_shareBuffer_sbuf_p0_rdat_950 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_951 = {_zz_shareBuffer_sbuf_p0_rdat_952,_zz_shareBuffer_sbuf_p0_rdat_953};
  assign _zz_shareBuffer_sbuf_p0_rdat_1063 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1064 = {_zz_shareBuffer_sbuf_p0_rdat_1065,_zz_shareBuffer_sbuf_p0_rdat_1066};
  assign _zz_shareBuffer_sbuf_p0_rdat_1177 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1178 = {_zz_shareBuffer_sbuf_p0_rdat_1179,_zz_shareBuffer_sbuf_p0_rdat_1180};
  assign _zz_shareBuffer_sbuf_p0_rdat_1290 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1291 = {_zz_shareBuffer_sbuf_p0_rdat_1292,_zz_shareBuffer_sbuf_p0_rdat_1293};
  assign _zz_shareBuffer_sbuf_p0_rdat_1403 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1404 = {_zz_shareBuffer_sbuf_p0_rdat_1405,_zz_shareBuffer_sbuf_p0_rdat_1406};
  assign _zz_shareBuffer_sbuf_p0_rdat_1515 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1516 = {_zz_shareBuffer_sbuf_p0_rdat_1517,_zz_shareBuffer_sbuf_p0_rdat_1518};
  assign _zz_shareBuffer_sbuf_p0_rdat_1627 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1628 = {_zz_shareBuffer_sbuf_p0_rdat_1629,_zz_shareBuffer_sbuf_p0_rdat_1630};
  assign _zz_shareBuffer_sbuf_p0_rdat_1737 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1738 = {_zz_shareBuffer_sbuf_p0_rdat_1739,_zz_shareBuffer_sbuf_p0_rdat_1740};
  assign _zz_shareBuffer_sbuf_p0_rdat_54 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_55 = {_zz_shareBuffer_sbuf_p0_rdat_56,_zz_shareBuffer_sbuf_p0_rdat_57};
  assign _zz_shareBuffer_sbuf_p0_rdat_163 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_164 = {_zz_shareBuffer_sbuf_p0_rdat_165,_zz_shareBuffer_sbuf_p0_rdat_166};
  assign _zz_shareBuffer_sbuf_p0_rdat_274 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_275 = {_zz_shareBuffer_sbuf_p0_rdat_276,_zz_shareBuffer_sbuf_p0_rdat_277};
  assign _zz_shareBuffer_sbuf_p0_rdat_385 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_386 = {_zz_shareBuffer_sbuf_p0_rdat_387,_zz_shareBuffer_sbuf_p0_rdat_388};
  assign _zz_shareBuffer_sbuf_p0_rdat_498 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_499 = {_zz_shareBuffer_sbuf_p0_rdat_500,_zz_shareBuffer_sbuf_p0_rdat_501};
  assign _zz_shareBuffer_sbuf_p0_rdat_611 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_612 = {_zz_shareBuffer_sbuf_p0_rdat_613,_zz_shareBuffer_sbuf_p0_rdat_614};
  assign _zz_shareBuffer_sbuf_p0_rdat_724 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_725 = {_zz_shareBuffer_sbuf_p0_rdat_726,_zz_shareBuffer_sbuf_p0_rdat_727};
  assign _zz_shareBuffer_sbuf_p0_rdat_837 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_838 = {_zz_shareBuffer_sbuf_p0_rdat_839,_zz_shareBuffer_sbuf_p0_rdat_840};
  assign _zz_shareBuffer_sbuf_p0_rdat_952 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_953 = {_zz_shareBuffer_sbuf_p0_rdat_954,_zz_shareBuffer_sbuf_p0_rdat_955};
  assign _zz_shareBuffer_sbuf_p0_rdat_1065 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1066 = {_zz_shareBuffer_sbuf_p0_rdat_1067,_zz_shareBuffer_sbuf_p0_rdat_1068};
  assign _zz_shareBuffer_sbuf_p0_rdat_1179 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1180 = {_zz_shareBuffer_sbuf_p0_rdat_1181,_zz_shareBuffer_sbuf_p0_rdat_1182};
  assign _zz_shareBuffer_sbuf_p0_rdat_1292 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1293 = {_zz_shareBuffer_sbuf_p0_rdat_1294,_zz_shareBuffer_sbuf_p0_rdat_1295};
  assign _zz_shareBuffer_sbuf_p0_rdat_1405 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1406 = {_zz_shareBuffer_sbuf_p0_rdat_1407,_zz_shareBuffer_sbuf_p0_rdat_1408};
  assign _zz_shareBuffer_sbuf_p0_rdat_1517 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1518 = {_zz_shareBuffer_sbuf_p0_rdat_1519,_zz_shareBuffer_sbuf_p0_rdat_1520};
  assign _zz_shareBuffer_sbuf_p0_rdat_1629 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1630 = {_zz_shareBuffer_sbuf_p0_rdat_1631,_zz_shareBuffer_sbuf_p0_rdat_1632};
  assign _zz_shareBuffer_sbuf_p0_rdat_1739 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1740 = {_zz_shareBuffer_sbuf_p0_rdat_1741,_zz_shareBuffer_sbuf_p0_rdat_1742};
  assign _zz_shareBuffer_sbuf_p0_rdat_56 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_57 = {_zz_shareBuffer_sbuf_p0_rdat_58,_zz_shareBuffer_sbuf_p0_rdat_59};
  assign _zz_shareBuffer_sbuf_p0_rdat_165 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_166 = {_zz_shareBuffer_sbuf_p0_rdat_167,_zz_shareBuffer_sbuf_p0_rdat_168};
  assign _zz_shareBuffer_sbuf_p0_rdat_276 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_277 = {_zz_shareBuffer_sbuf_p0_rdat_278,_zz_shareBuffer_sbuf_p0_rdat_279};
  assign _zz_shareBuffer_sbuf_p0_rdat_387 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_388 = {_zz_shareBuffer_sbuf_p0_rdat_389,_zz_shareBuffer_sbuf_p0_rdat_390};
  assign _zz_shareBuffer_sbuf_p0_rdat_500 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_501 = {_zz_shareBuffer_sbuf_p0_rdat_502,_zz_shareBuffer_sbuf_p0_rdat_503};
  assign _zz_shareBuffer_sbuf_p0_rdat_613 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_614 = {_zz_shareBuffer_sbuf_p0_rdat_615,_zz_shareBuffer_sbuf_p0_rdat_616};
  assign _zz_shareBuffer_sbuf_p0_rdat_726 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_727 = {_zz_shareBuffer_sbuf_p0_rdat_728,_zz_shareBuffer_sbuf_p0_rdat_729};
  assign _zz_shareBuffer_sbuf_p0_rdat_839 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_840 = {_zz_shareBuffer_sbuf_p0_rdat_841,_zz_shareBuffer_sbuf_p0_rdat_842};
  assign _zz_shareBuffer_sbuf_p0_rdat_954 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_955 = {_zz_shareBuffer_sbuf_p0_rdat_956,_zz_shareBuffer_sbuf_p0_rdat_957};
  assign _zz_shareBuffer_sbuf_p0_rdat_1067 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1068 = {_zz_shareBuffer_sbuf_p0_rdat_1069,_zz_shareBuffer_sbuf_p0_rdat_1070};
  assign _zz_shareBuffer_sbuf_p0_rdat_1181 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1182 = {_zz_shareBuffer_sbuf_p0_rdat_1183,_zz_shareBuffer_sbuf_p0_rdat_1184};
  assign _zz_shareBuffer_sbuf_p0_rdat_1294 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1295 = {_zz_shareBuffer_sbuf_p0_rdat_1296,_zz_shareBuffer_sbuf_p0_rdat_1297};
  assign _zz_shareBuffer_sbuf_p0_rdat_1407 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1408 = {_zz_shareBuffer_sbuf_p0_rdat_1409,_zz_shareBuffer_sbuf_p0_rdat_1410};
  assign _zz_shareBuffer_sbuf_p0_rdat_1519 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1520 = {_zz_shareBuffer_sbuf_p0_rdat_1521,_zz_shareBuffer_sbuf_p0_rdat_1522};
  assign _zz_shareBuffer_sbuf_p0_rdat_1631 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1632 = {_zz_shareBuffer_sbuf_p0_rdat_1633,_zz_shareBuffer_sbuf_p0_rdat_1634};
  assign _zz_shareBuffer_sbuf_p0_rdat_1741 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1742 = {_zz_shareBuffer_sbuf_p0_rdat_1743,_zz_shareBuffer_sbuf_p0_rdat_1744};
  assign _zz_shareBuffer_sbuf_p0_rdat_58 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_59 = {_zz_shareBuffer_sbuf_p0_rdat_60,_zz_shareBuffer_sbuf_p0_rdat_61};
  assign _zz_shareBuffer_sbuf_p0_rdat_167 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_168 = {_zz_shareBuffer_sbuf_p0_rdat_169,_zz_shareBuffer_sbuf_p0_rdat_170};
  assign _zz_shareBuffer_sbuf_p0_rdat_278 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_279 = {_zz_shareBuffer_sbuf_p0_rdat_280,_zz_shareBuffer_sbuf_p0_rdat_281};
  assign _zz_shareBuffer_sbuf_p0_rdat_389 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_390 = {_zz_shareBuffer_sbuf_p0_rdat_391,_zz_shareBuffer_sbuf_p0_rdat_392};
  assign _zz_shareBuffer_sbuf_p0_rdat_502 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_503 = {_zz_shareBuffer_sbuf_p0_rdat_504,_zz_shareBuffer_sbuf_p0_rdat_505};
  assign _zz_shareBuffer_sbuf_p0_rdat_615 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_616 = {_zz_shareBuffer_sbuf_p0_rdat_617,_zz_shareBuffer_sbuf_p0_rdat_618};
  assign _zz_shareBuffer_sbuf_p0_rdat_728 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_729 = {_zz_shareBuffer_sbuf_p0_rdat_730,_zz_shareBuffer_sbuf_p0_rdat_731};
  assign _zz_shareBuffer_sbuf_p0_rdat_841 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_842 = {_zz_shareBuffer_sbuf_p0_rdat_843,_zz_shareBuffer_sbuf_p0_rdat_844};
  assign _zz_shareBuffer_sbuf_p0_rdat_956 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_957 = {_zz_shareBuffer_sbuf_p0_rdat_958,_zz_shareBuffer_sbuf_p0_rdat_959};
  assign _zz_shareBuffer_sbuf_p0_rdat_1069 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1070 = {_zz_shareBuffer_sbuf_p0_rdat_1071,_zz_shareBuffer_sbuf_p0_rdat_1072};
  assign _zz_shareBuffer_sbuf_p0_rdat_1183 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1184 = {_zz_shareBuffer_sbuf_p0_rdat_1185,_zz_shareBuffer_sbuf_p0_rdat_1186};
  assign _zz_shareBuffer_sbuf_p0_rdat_1296 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1297 = {_zz_shareBuffer_sbuf_p0_rdat_1298,_zz_shareBuffer_sbuf_p0_rdat_1299};
  assign _zz_shareBuffer_sbuf_p0_rdat_1409 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1410 = {_zz_shareBuffer_sbuf_p0_rdat_1411,_zz_shareBuffer_sbuf_p0_rdat_1412};
  assign _zz_shareBuffer_sbuf_p0_rdat_1521 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1522 = {_zz_shareBuffer_sbuf_p0_rdat_1523,_zz_shareBuffer_sbuf_p0_rdat_1524};
  assign _zz_shareBuffer_sbuf_p0_rdat_1633 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1634 = {_zz_shareBuffer_sbuf_p0_rdat_1635,_zz_shareBuffer_sbuf_p0_rdat_1636};
  assign _zz_shareBuffer_sbuf_p0_rdat_1743 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1744 = {_zz_shareBuffer_sbuf_p0_rdat_1745,_zz_shareBuffer_sbuf_p0_rdat_1746};
  assign _zz_shareBuffer_sbuf_p0_rdat_60 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_61 = {_zz_shareBuffer_sbuf_p0_rdat_62,_zz_shareBuffer_sbuf_p0_rdat_63};
  assign _zz_shareBuffer_sbuf_p0_rdat_169 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_170 = {_zz_shareBuffer_sbuf_p0_rdat_171,_zz_shareBuffer_sbuf_p0_rdat_172};
  assign _zz_shareBuffer_sbuf_p0_rdat_280 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_281 = {_zz_shareBuffer_sbuf_p0_rdat_282,_zz_shareBuffer_sbuf_p0_rdat_283};
  assign _zz_shareBuffer_sbuf_p0_rdat_391 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_392 = {_zz_shareBuffer_sbuf_p0_rdat_393,_zz_shareBuffer_sbuf_p0_rdat_394};
  assign _zz_shareBuffer_sbuf_p0_rdat_504 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_505 = {_zz_shareBuffer_sbuf_p0_rdat_506,_zz_shareBuffer_sbuf_p0_rdat_507};
  assign _zz_shareBuffer_sbuf_p0_rdat_617 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_618 = {_zz_shareBuffer_sbuf_p0_rdat_619,_zz_shareBuffer_sbuf_p0_rdat_620};
  assign _zz_shareBuffer_sbuf_p0_rdat_730 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_731 = {_zz_shareBuffer_sbuf_p0_rdat_732,_zz_shareBuffer_sbuf_p0_rdat_733};
  assign _zz_shareBuffer_sbuf_p0_rdat_843 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_844 = {_zz_shareBuffer_sbuf_p0_rdat_845,_zz_shareBuffer_sbuf_p0_rdat_846};
  assign _zz_shareBuffer_sbuf_p0_rdat_958 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_959 = {_zz_shareBuffer_sbuf_p0_rdat_960,_zz_shareBuffer_sbuf_p0_rdat_961};
  assign _zz_shareBuffer_sbuf_p0_rdat_1071 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1072 = {_zz_shareBuffer_sbuf_p0_rdat_1073,_zz_shareBuffer_sbuf_p0_rdat_1074};
  assign _zz_shareBuffer_sbuf_p0_rdat_1185 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1186 = {_zz_shareBuffer_sbuf_p0_rdat_1187,_zz_shareBuffer_sbuf_p0_rdat_1188};
  assign _zz_shareBuffer_sbuf_p0_rdat_1298 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1299 = {_zz_shareBuffer_sbuf_p0_rdat_1300,_zz_shareBuffer_sbuf_p0_rdat_1301};
  assign _zz_shareBuffer_sbuf_p0_rdat_1411 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1412 = {_zz_shareBuffer_sbuf_p0_rdat_1413,_zz_shareBuffer_sbuf_p0_rdat_1414};
  assign _zz_shareBuffer_sbuf_p0_rdat_1523 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1524 = {_zz_shareBuffer_sbuf_p0_rdat_1525,_zz_shareBuffer_sbuf_p0_rdat_1526};
  assign _zz_shareBuffer_sbuf_p0_rdat_1635 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1636 = {_zz_shareBuffer_sbuf_p0_rdat_1637,_zz_shareBuffer_sbuf_p0_rdat_1638};
  assign _zz_shareBuffer_sbuf_p0_rdat_1745 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1746 = {_zz_shareBuffer_sbuf_p0_rdat_1747,_zz_shareBuffer_sbuf_p0_rdat_1748};
  assign _zz_shareBuffer_sbuf_p0_rdat_62 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_63 = {_zz_shareBuffer_sbuf_p0_rdat_64,_zz_shareBuffer_sbuf_p0_rdat_65};
  assign _zz_shareBuffer_sbuf_p0_rdat_171 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_172 = {_zz_shareBuffer_sbuf_p0_rdat_173,_zz_shareBuffer_sbuf_p0_rdat_174};
  assign _zz_shareBuffer_sbuf_p0_rdat_282 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_283 = {_zz_shareBuffer_sbuf_p0_rdat_284,_zz_shareBuffer_sbuf_p0_rdat_285};
  assign _zz_shareBuffer_sbuf_p0_rdat_393 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_394 = {_zz_shareBuffer_sbuf_p0_rdat_395,_zz_shareBuffer_sbuf_p0_rdat_396};
  assign _zz_shareBuffer_sbuf_p0_rdat_506 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_507 = {_zz_shareBuffer_sbuf_p0_rdat_508,_zz_shareBuffer_sbuf_p0_rdat_509};
  assign _zz_shareBuffer_sbuf_p0_rdat_619 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_620 = {_zz_shareBuffer_sbuf_p0_rdat_621,_zz_shareBuffer_sbuf_p0_rdat_622};
  assign _zz_shareBuffer_sbuf_p0_rdat_732 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_733 = {_zz_shareBuffer_sbuf_p0_rdat_734,_zz_shareBuffer_sbuf_p0_rdat_735};
  assign _zz_shareBuffer_sbuf_p0_rdat_845 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_846 = {_zz_shareBuffer_sbuf_p0_rdat_847,_zz_shareBuffer_sbuf_p0_rdat_848};
  assign _zz_shareBuffer_sbuf_p0_rdat_960 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_961 = {_zz_shareBuffer_sbuf_p0_rdat_962,_zz_shareBuffer_sbuf_p0_rdat_963};
  assign _zz_shareBuffer_sbuf_p0_rdat_1073 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1074 = {_zz_shareBuffer_sbuf_p0_rdat_1075,_zz_shareBuffer_sbuf_p0_rdat_1076};
  assign _zz_shareBuffer_sbuf_p0_rdat_1187 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1188 = {_zz_shareBuffer_sbuf_p0_rdat_1189,_zz_shareBuffer_sbuf_p0_rdat_1190};
  assign _zz_shareBuffer_sbuf_p0_rdat_1300 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1301 = {_zz_shareBuffer_sbuf_p0_rdat_1302,_zz_shareBuffer_sbuf_p0_rdat_1303};
  assign _zz_shareBuffer_sbuf_p0_rdat_1413 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1414 = {_zz_shareBuffer_sbuf_p0_rdat_1415,_zz_shareBuffer_sbuf_p0_rdat_1416};
  assign _zz_shareBuffer_sbuf_p0_rdat_1525 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1526 = {_zz_shareBuffer_sbuf_p0_rdat_1527,_zz_shareBuffer_sbuf_p0_rdat_1528};
  assign _zz_shareBuffer_sbuf_p0_rdat_1637 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1638 = {_zz_shareBuffer_sbuf_p0_rdat_1639,_zz_shareBuffer_sbuf_p0_rdat_1640};
  assign _zz_shareBuffer_sbuf_p0_rdat_1747 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1748 = {_zz_shareBuffer_sbuf_p0_rdat_1749,_zz_shareBuffer_sbuf_p0_rdat_1750};
  assign _zz_shareBuffer_sbuf_p0_rdat_64 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_65 = {_zz_shareBuffer_sbuf_p0_rdat_66,_zz_shareBuffer_sbuf_p0_rdat_67};
  assign _zz_shareBuffer_sbuf_p0_rdat_173 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_174 = {_zz_shareBuffer_sbuf_p0_rdat_175,_zz_shareBuffer_sbuf_p0_rdat_176};
  assign _zz_shareBuffer_sbuf_p0_rdat_284 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_285 = {_zz_shareBuffer_sbuf_p0_rdat_286,_zz_shareBuffer_sbuf_p0_rdat_287};
  assign _zz_shareBuffer_sbuf_p0_rdat_395 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_396 = {_zz_shareBuffer_sbuf_p0_rdat_397,_zz_shareBuffer_sbuf_p0_rdat_398};
  assign _zz_shareBuffer_sbuf_p0_rdat_508 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_509 = {_zz_shareBuffer_sbuf_p0_rdat_510,_zz_shareBuffer_sbuf_p0_rdat_511};
  assign _zz_shareBuffer_sbuf_p0_rdat_621 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_622 = {_zz_shareBuffer_sbuf_p0_rdat_623,_zz_shareBuffer_sbuf_p0_rdat_624};
  assign _zz_shareBuffer_sbuf_p0_rdat_734 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_735 = {_zz_shareBuffer_sbuf_p0_rdat_736,_zz_shareBuffer_sbuf_p0_rdat_737};
  assign _zz_shareBuffer_sbuf_p0_rdat_847 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_848 = {_zz_shareBuffer_sbuf_p0_rdat_849,_zz_shareBuffer_sbuf_p0_rdat_850};
  assign _zz_shareBuffer_sbuf_p0_rdat_962 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_963 = {_zz_shareBuffer_sbuf_p0_rdat_964,_zz_shareBuffer_sbuf_p0_rdat_965};
  assign _zz_shareBuffer_sbuf_p0_rdat_1075 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1076 = {_zz_shareBuffer_sbuf_p0_rdat_1077,_zz_shareBuffer_sbuf_p0_rdat_1078};
  assign _zz_shareBuffer_sbuf_p0_rdat_1189 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1190 = {_zz_shareBuffer_sbuf_p0_rdat_1191,_zz_shareBuffer_sbuf_p0_rdat_1192};
  assign _zz_shareBuffer_sbuf_p0_rdat_1302 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1303 = {_zz_shareBuffer_sbuf_p0_rdat_1304,_zz_shareBuffer_sbuf_p0_rdat_1305};
  assign _zz_shareBuffer_sbuf_p0_rdat_1415 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1416 = {_zz_shareBuffer_sbuf_p0_rdat_1417,_zz_shareBuffer_sbuf_p0_rdat_1418};
  assign _zz_shareBuffer_sbuf_p0_rdat_1527 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1528 = {_zz_shareBuffer_sbuf_p0_rdat_1529,_zz_shareBuffer_sbuf_p0_rdat_1530};
  assign _zz_shareBuffer_sbuf_p0_rdat_1639 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1640 = {_zz_shareBuffer_sbuf_p0_rdat_1641,_zz_shareBuffer_sbuf_p0_rdat_1642};
  assign _zz_shareBuffer_sbuf_p0_rdat_1749 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1750 = {_zz_shareBuffer_sbuf_p0_rdat_1751,_zz_shareBuffer_sbuf_p0_rdat_1752};
  assign _zz_shareBuffer_sbuf_p0_rdat_66 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_67 = {_zz_shareBuffer_sbuf_p0_rdat_68,_zz_shareBuffer_sbuf_p0_rdat_69};
  assign _zz_shareBuffer_sbuf_p0_rdat_175 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_176 = {_zz_shareBuffer_sbuf_p0_rdat_177,_zz_shareBuffer_sbuf_p0_rdat_178};
  assign _zz_shareBuffer_sbuf_p0_rdat_286 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_287 = {_zz_shareBuffer_sbuf_p0_rdat_288,_zz_shareBuffer_sbuf_p0_rdat_289};
  assign _zz_shareBuffer_sbuf_p0_rdat_397 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_398 = {_zz_shareBuffer_sbuf_p0_rdat_399,_zz_shareBuffer_sbuf_p0_rdat_400};
  assign _zz_shareBuffer_sbuf_p0_rdat_510 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_511 = {_zz_shareBuffer_sbuf_p0_rdat_512,_zz_shareBuffer_sbuf_p0_rdat_513};
  assign _zz_shareBuffer_sbuf_p0_rdat_623 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_624 = {_zz_shareBuffer_sbuf_p0_rdat_625,_zz_shareBuffer_sbuf_p0_rdat_626};
  assign _zz_shareBuffer_sbuf_p0_rdat_736 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_737 = {_zz_shareBuffer_sbuf_p0_rdat_738,_zz_shareBuffer_sbuf_p0_rdat_739};
  assign _zz_shareBuffer_sbuf_p0_rdat_849 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_850 = {_zz_shareBuffer_sbuf_p0_rdat_851,_zz_shareBuffer_sbuf_p0_rdat_852};
  assign _zz_shareBuffer_sbuf_p0_rdat_964 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_965 = {_zz_shareBuffer_sbuf_p0_rdat_966,_zz_shareBuffer_sbuf_p0_rdat_967};
  assign _zz_shareBuffer_sbuf_p0_rdat_1077 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1078 = {_zz_shareBuffer_sbuf_p0_rdat_1079,_zz_shareBuffer_sbuf_p0_rdat_1080};
  assign _zz_shareBuffer_sbuf_p0_rdat_1191 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1192 = {_zz_shareBuffer_sbuf_p0_rdat_1193,_zz_shareBuffer_sbuf_p0_rdat_1194};
  assign _zz_shareBuffer_sbuf_p0_rdat_1304 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1305 = {_zz_shareBuffer_sbuf_p0_rdat_1306,_zz_shareBuffer_sbuf_p0_rdat_1307};
  assign _zz_shareBuffer_sbuf_p0_rdat_1417 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1418 = {_zz_shareBuffer_sbuf_p0_rdat_1419,_zz_shareBuffer_sbuf_p0_rdat_1420};
  assign _zz_shareBuffer_sbuf_p0_rdat_1529 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1530 = {_zz_shareBuffer_sbuf_p0_rdat_1531,_zz_shareBuffer_sbuf_p0_rdat_1532};
  assign _zz_shareBuffer_sbuf_p0_rdat_1641 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1642 = {_zz_shareBuffer_sbuf_p0_rdat_1643,_zz_shareBuffer_sbuf_p0_rdat_1644};
  assign _zz_shareBuffer_sbuf_p0_rdat_1751 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1752 = {_zz_shareBuffer_sbuf_p0_rdat_1753,_zz_shareBuffer_sbuf_p0_rdat_1754};
  assign _zz_shareBuffer_sbuf_p0_rdat_68 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_69 = {_zz_shareBuffer_sbuf_p0_rdat_70,_zz_shareBuffer_sbuf_p0_rdat_71};
  assign _zz_shareBuffer_sbuf_p0_rdat_177 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_178 = {_zz_shareBuffer_sbuf_p0_rdat_179,_zz_shareBuffer_sbuf_p0_rdat_180};
  assign _zz_shareBuffer_sbuf_p0_rdat_288 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_289 = {_zz_shareBuffer_sbuf_p0_rdat_290,_zz_shareBuffer_sbuf_p0_rdat_291};
  assign _zz_shareBuffer_sbuf_p0_rdat_399 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_400 = {_zz_shareBuffer_sbuf_p0_rdat_401,_zz_shareBuffer_sbuf_p0_rdat_402};
  assign _zz_shareBuffer_sbuf_p0_rdat_512 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_513 = {_zz_shareBuffer_sbuf_p0_rdat_514,_zz_shareBuffer_sbuf_p0_rdat_515};
  assign _zz_shareBuffer_sbuf_p0_rdat_625 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_626 = {_zz_shareBuffer_sbuf_p0_rdat_627,_zz_shareBuffer_sbuf_p0_rdat_628};
  assign _zz_shareBuffer_sbuf_p0_rdat_738 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_739 = {_zz_shareBuffer_sbuf_p0_rdat_740,_zz_shareBuffer_sbuf_p0_rdat_741};
  assign _zz_shareBuffer_sbuf_p0_rdat_851 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_852 = {_zz_shareBuffer_sbuf_p0_rdat_853,_zz_shareBuffer_sbuf_p0_rdat_854};
  assign _zz_shareBuffer_sbuf_p0_rdat_966 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_967 = {_zz_shareBuffer_sbuf_p0_rdat_968,_zz_shareBuffer_sbuf_p0_rdat_969};
  assign _zz_shareBuffer_sbuf_p0_rdat_1079 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1080 = {_zz_shareBuffer_sbuf_p0_rdat_1081,_zz_shareBuffer_sbuf_p0_rdat_1082};
  assign _zz_shareBuffer_sbuf_p0_rdat_1193 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1194 = {_zz_shareBuffer_sbuf_p0_rdat_1195,_zz_shareBuffer_sbuf_p0_rdat_1196};
  assign _zz_shareBuffer_sbuf_p0_rdat_1306 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1307 = {_zz_shareBuffer_sbuf_p0_rdat_1308,_zz_shareBuffer_sbuf_p0_rdat_1309};
  assign _zz_shareBuffer_sbuf_p0_rdat_1419 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1420 = {_zz_shareBuffer_sbuf_p0_rdat_1421,_zz_shareBuffer_sbuf_p0_rdat_1422};
  assign _zz_shareBuffer_sbuf_p0_rdat_1531 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1532 = {_zz_shareBuffer_sbuf_p0_rdat_1533,_zz_shareBuffer_sbuf_p0_rdat_1534};
  assign _zz_shareBuffer_sbuf_p0_rdat_1643 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1644 = {_zz_shareBuffer_sbuf_p0_rdat_1645,_zz_shareBuffer_sbuf_p0_rdat_1646};
  assign _zz_shareBuffer_sbuf_p0_rdat_1753 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1754 = {_zz_shareBuffer_sbuf_p0_rdat_1755,_zz_shareBuffer_sbuf_p0_rdat_1756};
  assign _zz_shareBuffer_sbuf_p0_rdat_70 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_71 = {_zz_shareBuffer_sbuf_p0_rdat_72,_zz_shareBuffer_sbuf_p0_rdat_73};
  assign _zz_shareBuffer_sbuf_p0_rdat_179 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_180 = {_zz_shareBuffer_sbuf_p0_rdat_181,_zz_shareBuffer_sbuf_p0_rdat_182};
  assign _zz_shareBuffer_sbuf_p0_rdat_290 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_291 = {_zz_shareBuffer_sbuf_p0_rdat_292,_zz_shareBuffer_sbuf_p0_rdat_293};
  assign _zz_shareBuffer_sbuf_p0_rdat_401 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_402 = {_zz_shareBuffer_sbuf_p0_rdat_403,_zz_shareBuffer_sbuf_p0_rdat_404};
  assign _zz_shareBuffer_sbuf_p0_rdat_514 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_515 = {_zz_shareBuffer_sbuf_p0_rdat_516,_zz_shareBuffer_sbuf_p0_rdat_517};
  assign _zz_shareBuffer_sbuf_p0_rdat_627 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_628 = {_zz_shareBuffer_sbuf_p0_rdat_629,_zz_shareBuffer_sbuf_p0_rdat_630};
  assign _zz_shareBuffer_sbuf_p0_rdat_740 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_741 = {_zz_shareBuffer_sbuf_p0_rdat_742,_zz_shareBuffer_sbuf_p0_rdat_743};
  assign _zz_shareBuffer_sbuf_p0_rdat_853 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_854 = {_zz_shareBuffer_sbuf_p0_rdat_855,_zz_shareBuffer_sbuf_p0_rdat_856};
  assign _zz_shareBuffer_sbuf_p0_rdat_968 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_969 = {_zz_shareBuffer_sbuf_p0_rdat_970,_zz_shareBuffer_sbuf_p0_rdat_971};
  assign _zz_shareBuffer_sbuf_p0_rdat_1081 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1082 = {_zz_shareBuffer_sbuf_p0_rdat_1083,_zz_shareBuffer_sbuf_p0_rdat_1084};
  assign _zz_shareBuffer_sbuf_p0_rdat_1195 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1196 = {_zz_shareBuffer_sbuf_p0_rdat_1197,_zz_shareBuffer_sbuf_p0_rdat_1198};
  assign _zz_shareBuffer_sbuf_p0_rdat_1308 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1309 = {_zz_shareBuffer_sbuf_p0_rdat_1310,_zz_shareBuffer_sbuf_p0_rdat_1311};
  assign _zz_shareBuffer_sbuf_p0_rdat_1421 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1422 = {_zz_shareBuffer_sbuf_p0_rdat_1423,_zz_shareBuffer_sbuf_p0_rdat_1424};
  assign _zz_shareBuffer_sbuf_p0_rdat_1533 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1534 = {_zz_shareBuffer_sbuf_p0_rdat_1535,_zz_shareBuffer_sbuf_p0_rdat_1536};
  assign _zz_shareBuffer_sbuf_p0_rdat_1645 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1646 = {_zz_shareBuffer_sbuf_p0_rdat_1647,_zz_shareBuffer_sbuf_p0_rdat_1648};
  assign _zz_shareBuffer_sbuf_p0_rdat_1755 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1756 = {_zz_shareBuffer_sbuf_p0_rdat_1757,_zz_shareBuffer_sbuf_p0_rdat_1758};
  assign _zz_shareBuffer_sbuf_p0_rdat_72 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_73 = {_zz_shareBuffer_sbuf_p0_rdat_74,_zz_shareBuffer_sbuf_p0_rdat_75};
  assign _zz_shareBuffer_sbuf_p0_rdat_181 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_182 = {_zz_shareBuffer_sbuf_p0_rdat_183,_zz_shareBuffer_sbuf_p0_rdat_184};
  assign _zz_shareBuffer_sbuf_p0_rdat_292 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_293 = {_zz_shareBuffer_sbuf_p0_rdat_294,_zz_shareBuffer_sbuf_p0_rdat_295};
  assign _zz_shareBuffer_sbuf_p0_rdat_403 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_404 = {_zz_shareBuffer_sbuf_p0_rdat_405,_zz_shareBuffer_sbuf_p0_rdat_406};
  assign _zz_shareBuffer_sbuf_p0_rdat_516 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_517 = {_zz_shareBuffer_sbuf_p0_rdat_518,_zz_shareBuffer_sbuf_p0_rdat_519};
  assign _zz_shareBuffer_sbuf_p0_rdat_629 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_630 = {_zz_shareBuffer_sbuf_p0_rdat_631,_zz_shareBuffer_sbuf_p0_rdat_632};
  assign _zz_shareBuffer_sbuf_p0_rdat_742 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_743 = {_zz_shareBuffer_sbuf_p0_rdat_744,_zz_shareBuffer_sbuf_p0_rdat_745};
  assign _zz_shareBuffer_sbuf_p0_rdat_855 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_856 = {_zz_shareBuffer_sbuf_p0_rdat_857,_zz_shareBuffer_sbuf_p0_rdat_858};
  assign _zz_shareBuffer_sbuf_p0_rdat_970 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_971 = {_zz_shareBuffer_sbuf_p0_rdat_972,_zz_shareBuffer_sbuf_p0_rdat_973};
  assign _zz_shareBuffer_sbuf_p0_rdat_1083 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1084 = {_zz_shareBuffer_sbuf_p0_rdat_1085,_zz_shareBuffer_sbuf_p0_rdat_1086};
  assign _zz_shareBuffer_sbuf_p0_rdat_1197 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1198 = {_zz_shareBuffer_sbuf_p0_rdat_1199,_zz_shareBuffer_sbuf_p0_rdat_1200};
  assign _zz_shareBuffer_sbuf_p0_rdat_1310 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1311 = {_zz_shareBuffer_sbuf_p0_rdat_1312,_zz_shareBuffer_sbuf_p0_rdat_1313};
  assign _zz_shareBuffer_sbuf_p0_rdat_1423 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1424 = {_zz_shareBuffer_sbuf_p0_rdat_1425,_zz_shareBuffer_sbuf_p0_rdat_1426};
  assign _zz_shareBuffer_sbuf_p0_rdat_1535 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1536 = {_zz_shareBuffer_sbuf_p0_rdat_1537,_zz_shareBuffer_sbuf_p0_rdat_1538};
  assign _zz_shareBuffer_sbuf_p0_rdat_1647 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1648 = {_zz_shareBuffer_sbuf_p0_rdat_1649,_zz_shareBuffer_sbuf_p0_rdat_1650};
  assign _zz_shareBuffer_sbuf_p0_rdat_1757 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1758 = {_zz_shareBuffer_sbuf_p0_rdat_1759,_zz_shareBuffer_sbuf_p0_rdat_1760};
  assign _zz_shareBuffer_sbuf_p0_rdat_74 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_75 = {_zz_shareBuffer_sbuf_p0_rdat_76,_zz_shareBuffer_sbuf_p0_rdat_77};
  assign _zz_shareBuffer_sbuf_p0_rdat_183 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_184 = {_zz_shareBuffer_sbuf_p0_rdat_185,_zz_shareBuffer_sbuf_p0_rdat_186};
  assign _zz_shareBuffer_sbuf_p0_rdat_294 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_295 = {_zz_shareBuffer_sbuf_p0_rdat_296,_zz_shareBuffer_sbuf_p0_rdat_297};
  assign _zz_shareBuffer_sbuf_p0_rdat_405 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_406 = {_zz_shareBuffer_sbuf_p0_rdat_407,_zz_shareBuffer_sbuf_p0_rdat_408};
  assign _zz_shareBuffer_sbuf_p0_rdat_518 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_519 = {_zz_shareBuffer_sbuf_p0_rdat_520,_zz_shareBuffer_sbuf_p0_rdat_521};
  assign _zz_shareBuffer_sbuf_p0_rdat_631 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_632 = {_zz_shareBuffer_sbuf_p0_rdat_633,_zz_shareBuffer_sbuf_p0_rdat_634};
  assign _zz_shareBuffer_sbuf_p0_rdat_744 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_745 = {_zz_shareBuffer_sbuf_p0_rdat_746,_zz_shareBuffer_sbuf_p0_rdat_747};
  assign _zz_shareBuffer_sbuf_p0_rdat_857 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_858 = {_zz_shareBuffer_sbuf_p0_rdat_859,_zz_shareBuffer_sbuf_p0_rdat_860};
  assign _zz_shareBuffer_sbuf_p0_rdat_972 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_973 = {_zz_shareBuffer_sbuf_p0_rdat_974,_zz_shareBuffer_sbuf_p0_rdat_975};
  assign _zz_shareBuffer_sbuf_p0_rdat_1085 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1086 = {_zz_shareBuffer_sbuf_p0_rdat_1087,_zz_shareBuffer_sbuf_p0_rdat_1088};
  assign _zz_shareBuffer_sbuf_p0_rdat_1199 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1200 = {_zz_shareBuffer_sbuf_p0_rdat_1201,_zz_shareBuffer_sbuf_p0_rdat_1202};
  assign _zz_shareBuffer_sbuf_p0_rdat_1312 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1313 = {_zz_shareBuffer_sbuf_p0_rdat_1314,_zz_shareBuffer_sbuf_p0_rdat_1315};
  assign _zz_shareBuffer_sbuf_p0_rdat_1425 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1426 = {_zz_shareBuffer_sbuf_p0_rdat_1427,_zz_shareBuffer_sbuf_p0_rdat_1428};
  assign _zz_shareBuffer_sbuf_p0_rdat_1537 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1538 = {_zz_shareBuffer_sbuf_p0_rdat_1539,_zz_shareBuffer_sbuf_p0_rdat_1540};
  assign _zz_shareBuffer_sbuf_p0_rdat_1649 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1650 = {_zz_shareBuffer_sbuf_p0_rdat_1651,_zz_shareBuffer_sbuf_p0_rdat_1652};
  assign _zz_shareBuffer_sbuf_p0_rdat_1759 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1760 = {_zz_shareBuffer_sbuf_p0_rdat_1761,_zz_shareBuffer_sbuf_p0_rdat_1762};
  assign _zz_shareBuffer_sbuf_p0_rdat_76 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_77 = {_zz_shareBuffer_sbuf_p0_rdat_78,_zz_shareBuffer_sbuf_p0_rdat_79};
  assign _zz_shareBuffer_sbuf_p0_rdat_185 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_186 = {_zz_shareBuffer_sbuf_p0_rdat_187,_zz_shareBuffer_sbuf_p0_rdat_188};
  assign _zz_shareBuffer_sbuf_p0_rdat_296 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_297 = {_zz_shareBuffer_sbuf_p0_rdat_298,_zz_shareBuffer_sbuf_p0_rdat_299};
  assign _zz_shareBuffer_sbuf_p0_rdat_407 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_408 = {_zz_shareBuffer_sbuf_p0_rdat_409,_zz_shareBuffer_sbuf_p0_rdat_410};
  assign _zz_shareBuffer_sbuf_p0_rdat_520 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_521 = {_zz_shareBuffer_sbuf_p0_rdat_522,_zz_shareBuffer_sbuf_p0_rdat_523};
  assign _zz_shareBuffer_sbuf_p0_rdat_633 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_634 = {_zz_shareBuffer_sbuf_p0_rdat_635,_zz_shareBuffer_sbuf_p0_rdat_636};
  assign _zz_shareBuffer_sbuf_p0_rdat_746 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_747 = {_zz_shareBuffer_sbuf_p0_rdat_748,_zz_shareBuffer_sbuf_p0_rdat_749};
  assign _zz_shareBuffer_sbuf_p0_rdat_859 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_860 = {_zz_shareBuffer_sbuf_p0_rdat_861,_zz_shareBuffer_sbuf_p0_rdat_862};
  assign _zz_shareBuffer_sbuf_p0_rdat_974 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_975 = {_zz_shareBuffer_sbuf_p0_rdat_976,_zz_shareBuffer_sbuf_p0_rdat_977};
  assign _zz_shareBuffer_sbuf_p0_rdat_1087 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1088 = {_zz_shareBuffer_sbuf_p0_rdat_1089,_zz_shareBuffer_sbuf_p0_rdat_1090};
  assign _zz_shareBuffer_sbuf_p0_rdat_1201 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1202 = {_zz_shareBuffer_sbuf_p0_rdat_1203,_zz_shareBuffer_sbuf_p0_rdat_1204};
  assign _zz_shareBuffer_sbuf_p0_rdat_1314 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1315 = {_zz_shareBuffer_sbuf_p0_rdat_1316,_zz_shareBuffer_sbuf_p0_rdat_1317};
  assign _zz_shareBuffer_sbuf_p0_rdat_1427 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1428 = {_zz_shareBuffer_sbuf_p0_rdat_1429,_zz_shareBuffer_sbuf_p0_rdat_1430};
  assign _zz_shareBuffer_sbuf_p0_rdat_1539 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1540 = {_zz_shareBuffer_sbuf_p0_rdat_1541,_zz_shareBuffer_sbuf_p0_rdat_1542};
  assign _zz_shareBuffer_sbuf_p0_rdat_1651 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1652 = {_zz_shareBuffer_sbuf_p0_rdat_1653,_zz_shareBuffer_sbuf_p0_rdat_1654};
  assign _zz_shareBuffer_sbuf_p0_rdat_1761 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1762 = {_zz_shareBuffer_sbuf_p0_rdat_1763,_zz_shareBuffer_sbuf_p0_rdat_1764};
  assign _zz_shareBuffer_sbuf_p0_rdat_78 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_79 = {_zz_shareBuffer_sbuf_p0_rdat_80,_zz_shareBuffer_sbuf_p0_rdat_81};
  assign _zz_shareBuffer_sbuf_p0_rdat_187 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_188 = {_zz_shareBuffer_sbuf_p0_rdat_189,_zz_shareBuffer_sbuf_p0_rdat_190};
  assign _zz_shareBuffer_sbuf_p0_rdat_298 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_299 = {_zz_shareBuffer_sbuf_p0_rdat_300,_zz_shareBuffer_sbuf_p0_rdat_301};
  assign _zz_shareBuffer_sbuf_p0_rdat_409 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_410 = {_zz_shareBuffer_sbuf_p0_rdat_411,_zz_shareBuffer_sbuf_p0_rdat_412};
  assign _zz_shareBuffer_sbuf_p0_rdat_522 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_523 = {_zz_shareBuffer_sbuf_p0_rdat_524,_zz_shareBuffer_sbuf_p0_rdat_525};
  assign _zz_shareBuffer_sbuf_p0_rdat_635 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_636 = {_zz_shareBuffer_sbuf_p0_rdat_637,_zz_shareBuffer_sbuf_p0_rdat_638};
  assign _zz_shareBuffer_sbuf_p0_rdat_748 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_749 = {_zz_shareBuffer_sbuf_p0_rdat_750,_zz_shareBuffer_sbuf_p0_rdat_751};
  assign _zz_shareBuffer_sbuf_p0_rdat_861 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_862 = {_zz_shareBuffer_sbuf_p0_rdat_863,_zz_shareBuffer_sbuf_p0_rdat_864};
  assign _zz_shareBuffer_sbuf_p0_rdat_976 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_977 = {_zz_shareBuffer_sbuf_p0_rdat_978,_zz_shareBuffer_sbuf_p0_rdat_979};
  assign _zz_shareBuffer_sbuf_p0_rdat_1089 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1090 = {_zz_shareBuffer_sbuf_p0_rdat_1091,_zz_shareBuffer_sbuf_p0_rdat_1092};
  assign _zz_shareBuffer_sbuf_p0_rdat_1203 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1204 = {_zz_shareBuffer_sbuf_p0_rdat_1205,_zz_shareBuffer_sbuf_p0_rdat_1206};
  assign _zz_shareBuffer_sbuf_p0_rdat_1316 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1317 = {_zz_shareBuffer_sbuf_p0_rdat_1318,_zz_shareBuffer_sbuf_p0_rdat_1319};
  assign _zz_shareBuffer_sbuf_p0_rdat_1429 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1430 = {_zz_shareBuffer_sbuf_p0_rdat_1431,_zz_shareBuffer_sbuf_p0_rdat_1432};
  assign _zz_shareBuffer_sbuf_p0_rdat_1541 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1542 = {_zz_shareBuffer_sbuf_p0_rdat_1543,_zz_shareBuffer_sbuf_p0_rdat_1544};
  assign _zz_shareBuffer_sbuf_p0_rdat_1653 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1654 = {_zz_shareBuffer_sbuf_p0_rdat_1655,_zz_shareBuffer_sbuf_p0_rdat_1656};
  assign _zz_shareBuffer_sbuf_p0_rdat_1763 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1764 = {_zz_shareBuffer_sbuf_p0_rdat_1765,_zz_shareBuffer_sbuf_p0_rdat_1766};
  assign _zz_shareBuffer_sbuf_p0_rdat_80 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_81 = {_zz_shareBuffer_sbuf_p0_rdat_82,_zz_shareBuffer_sbuf_p0_rdat_83};
  assign _zz_shareBuffer_sbuf_p0_rdat_189 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_190 = {_zz_shareBuffer_sbuf_p0_rdat_191,_zz_shareBuffer_sbuf_p0_rdat_192};
  assign _zz_shareBuffer_sbuf_p0_rdat_300 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_301 = {_zz_shareBuffer_sbuf_p0_rdat_302,_zz_shareBuffer_sbuf_p0_rdat_303};
  assign _zz_shareBuffer_sbuf_p0_rdat_411 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_412 = {_zz_shareBuffer_sbuf_p0_rdat_413,_zz_shareBuffer_sbuf_p0_rdat_414};
  assign _zz_shareBuffer_sbuf_p0_rdat_524 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_525 = {_zz_shareBuffer_sbuf_p0_rdat_526,_zz_shareBuffer_sbuf_p0_rdat_527};
  assign _zz_shareBuffer_sbuf_p0_rdat_637 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_638 = {_zz_shareBuffer_sbuf_p0_rdat_639,_zz_shareBuffer_sbuf_p0_rdat_640};
  assign _zz_shareBuffer_sbuf_p0_rdat_750 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_751 = {_zz_shareBuffer_sbuf_p0_rdat_752,_zz_shareBuffer_sbuf_p0_rdat_753};
  assign _zz_shareBuffer_sbuf_p0_rdat_863 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_864 = {_zz_shareBuffer_sbuf_p0_rdat_865,_zz_shareBuffer_sbuf_p0_rdat_866};
  assign _zz_shareBuffer_sbuf_p0_rdat_978 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_979 = {_zz_shareBuffer_sbuf_p0_rdat_980,_zz_shareBuffer_sbuf_p0_rdat_981};
  assign _zz_shareBuffer_sbuf_p0_rdat_1091 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1092 = {_zz_shareBuffer_sbuf_p0_rdat_1093,_zz_shareBuffer_sbuf_p0_rdat_1094};
  assign _zz_shareBuffer_sbuf_p0_rdat_1205 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1206 = {_zz_shareBuffer_sbuf_p0_rdat_1207,_zz_shareBuffer_sbuf_p0_rdat_1208};
  assign _zz_shareBuffer_sbuf_p0_rdat_1318 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1319 = {_zz_shareBuffer_sbuf_p0_rdat_1320,_zz_shareBuffer_sbuf_p0_rdat_1321};
  assign _zz_shareBuffer_sbuf_p0_rdat_1431 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1432 = {_zz_shareBuffer_sbuf_p0_rdat_1433,_zz_shareBuffer_sbuf_p0_rdat_1434};
  assign _zz_shareBuffer_sbuf_p0_rdat_1543 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1544 = {_zz_shareBuffer_sbuf_p0_rdat_1545,_zz_shareBuffer_sbuf_p0_rdat_1546};
  assign _zz_shareBuffer_sbuf_p0_rdat_1655 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1656 = {_zz_shareBuffer_sbuf_p0_rdat_1657,_zz_shareBuffer_sbuf_p0_rdat_1658};
  assign _zz_shareBuffer_sbuf_p0_rdat_1765 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1766 = {_zz_shareBuffer_sbuf_p0_rdat_1767,_zz_shareBuffer_sbuf_p0_rdat_1768};
  assign _zz_shareBuffer_sbuf_p0_rdat_82 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_83 = {_zz_shareBuffer_sbuf_p0_rdat_84,_zz_shareBuffer_sbuf_p0_rdat_85};
  assign _zz_shareBuffer_sbuf_p0_rdat_191 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_192 = {_zz_shareBuffer_sbuf_p0_rdat_193,_zz_shareBuffer_sbuf_p0_rdat_194};
  assign _zz_shareBuffer_sbuf_p0_rdat_302 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_303 = {_zz_shareBuffer_sbuf_p0_rdat_304,_zz_shareBuffer_sbuf_p0_rdat_305};
  assign _zz_shareBuffer_sbuf_p0_rdat_413 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_414 = {_zz_shareBuffer_sbuf_p0_rdat_415,_zz_shareBuffer_sbuf_p0_rdat_416};
  assign _zz_shareBuffer_sbuf_p0_rdat_526 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_527 = {_zz_shareBuffer_sbuf_p0_rdat_528,_zz_shareBuffer_sbuf_p0_rdat_529};
  assign _zz_shareBuffer_sbuf_p0_rdat_639 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_640 = {_zz_shareBuffer_sbuf_p0_rdat_641,_zz_shareBuffer_sbuf_p0_rdat_642};
  assign _zz_shareBuffer_sbuf_p0_rdat_752 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_753 = {_zz_shareBuffer_sbuf_p0_rdat_754,_zz_shareBuffer_sbuf_p0_rdat_755};
  assign _zz_shareBuffer_sbuf_p0_rdat_865 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_866 = {_zz_shareBuffer_sbuf_p0_rdat_867,_zz_shareBuffer_sbuf_p0_rdat_868};
  assign _zz_shareBuffer_sbuf_p0_rdat_980 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_981 = {_zz_shareBuffer_sbuf_p0_rdat_982,_zz_shareBuffer_sbuf_p0_rdat_983};
  assign _zz_shareBuffer_sbuf_p0_rdat_1093 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1094 = {_zz_shareBuffer_sbuf_p0_rdat_1095,_zz_shareBuffer_sbuf_p0_rdat_1096};
  assign _zz_shareBuffer_sbuf_p0_rdat_1207 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1208 = {_zz_shareBuffer_sbuf_p0_rdat_1209,_zz_shareBuffer_sbuf_p0_rdat_1210};
  assign _zz_shareBuffer_sbuf_p0_rdat_1320 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1321 = {_zz_shareBuffer_sbuf_p0_rdat_1322,_zz_shareBuffer_sbuf_p0_rdat_1323};
  assign _zz_shareBuffer_sbuf_p0_rdat_1433 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1434 = {_zz_shareBuffer_sbuf_p0_rdat_1435,_zz_shareBuffer_sbuf_p0_rdat_1436};
  assign _zz_shareBuffer_sbuf_p0_rdat_1545 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1546 = {_zz_shareBuffer_sbuf_p0_rdat_1547,_zz_shareBuffer_sbuf_p0_rdat_1548};
  assign _zz_shareBuffer_sbuf_p0_rdat_1657 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1658 = {_zz_shareBuffer_sbuf_p0_rdat_1659,_zz_shareBuffer_sbuf_p0_rdat_1660};
  assign _zz_shareBuffer_sbuf_p0_rdat_1767 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1768 = {_zz_shareBuffer_sbuf_p0_rdat_1769,_zz_shareBuffer_sbuf_p0_rdat_1770};
  assign _zz_shareBuffer_sbuf_p0_rdat_84 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_85 = {_zz_shareBuffer_sbuf_p0_rdat_86,_zz_shareBuffer_sbuf_p0_rdat_87};
  assign _zz_shareBuffer_sbuf_p0_rdat_193 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_194 = {_zz_shareBuffer_sbuf_p0_rdat_195,_zz_shareBuffer_sbuf_p0_rdat_196};
  assign _zz_shareBuffer_sbuf_p0_rdat_304 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_305 = {_zz_shareBuffer_sbuf_p0_rdat_306,_zz_shareBuffer_sbuf_p0_rdat_307};
  assign _zz_shareBuffer_sbuf_p0_rdat_415 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_416 = {_zz_shareBuffer_sbuf_p0_rdat_417,_zz_shareBuffer_sbuf_p0_rdat_418};
  assign _zz_shareBuffer_sbuf_p0_rdat_528 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_529 = {_zz_shareBuffer_sbuf_p0_rdat_530,_zz_shareBuffer_sbuf_p0_rdat_531};
  assign _zz_shareBuffer_sbuf_p0_rdat_641 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_642 = {_zz_shareBuffer_sbuf_p0_rdat_643,_zz_shareBuffer_sbuf_p0_rdat_644};
  assign _zz_shareBuffer_sbuf_p0_rdat_754 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_755 = {_zz_shareBuffer_sbuf_p0_rdat_756,_zz_shareBuffer_sbuf_p0_rdat_757};
  assign _zz_shareBuffer_sbuf_p0_rdat_867 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_868 = {_zz_shareBuffer_sbuf_p0_rdat_869,_zz_shareBuffer_sbuf_p0_rdat_870};
  assign _zz_shareBuffer_sbuf_p0_rdat_982 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_983 = {_zz_shareBuffer_sbuf_p0_rdat_984,_zz_shareBuffer_sbuf_p0_rdat_985};
  assign _zz_shareBuffer_sbuf_p0_rdat_1095 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1096 = {_zz_shareBuffer_sbuf_p0_rdat_1097,_zz_shareBuffer_sbuf_p0_rdat_1098};
  assign _zz_shareBuffer_sbuf_p0_rdat_1209 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1210 = {_zz_shareBuffer_sbuf_p0_rdat_1211,_zz_shareBuffer_sbuf_p0_rdat_1212};
  assign _zz_shareBuffer_sbuf_p0_rdat_1322 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1323 = {_zz_shareBuffer_sbuf_p0_rdat_1324,_zz_shareBuffer_sbuf_p0_rdat_1325};
  assign _zz_shareBuffer_sbuf_p0_rdat_1435 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1436 = {_zz_shareBuffer_sbuf_p0_rdat_1437,_zz_shareBuffer_sbuf_p0_rdat_1438};
  assign _zz_shareBuffer_sbuf_p0_rdat_1547 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1548 = {_zz_shareBuffer_sbuf_p0_rdat_1549,_zz_shareBuffer_sbuf_p0_rdat_1550};
  assign _zz_shareBuffer_sbuf_p0_rdat_1659 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1660 = {_zz_shareBuffer_sbuf_p0_rdat_1661,_zz_shareBuffer_sbuf_p0_rdat_1662};
  assign _zz_shareBuffer_sbuf_p0_rdat_1769 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1770 = {_zz_shareBuffer_sbuf_p0_rdat_1771,_zz_shareBuffer_sbuf_p0_rdat_1772};
  assign _zz_shareBuffer_sbuf_p0_rdat_86 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_87 = {_zz_shareBuffer_sbuf_p0_rdat_88,_zz_shareBuffer_sbuf_p0_rdat_89};
  assign _zz_shareBuffer_sbuf_p0_rdat_195 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_196 = {_zz_shareBuffer_sbuf_p0_rdat_197,_zz_shareBuffer_sbuf_p0_rdat_198};
  assign _zz_shareBuffer_sbuf_p0_rdat_306 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_307 = {_zz_shareBuffer_sbuf_p0_rdat_308,_zz_shareBuffer_sbuf_p0_rdat_309};
  assign _zz_shareBuffer_sbuf_p0_rdat_417 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_418 = {_zz_shareBuffer_sbuf_p0_rdat_419,_zz_shareBuffer_sbuf_p0_rdat_420};
  assign _zz_shareBuffer_sbuf_p0_rdat_530 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_531 = {_zz_shareBuffer_sbuf_p0_rdat_532,_zz_shareBuffer_sbuf_p0_rdat_533};
  assign _zz_shareBuffer_sbuf_p0_rdat_643 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_644 = {_zz_shareBuffer_sbuf_p0_rdat_645,_zz_shareBuffer_sbuf_p0_rdat_646};
  assign _zz_shareBuffer_sbuf_p0_rdat_756 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_757 = {_zz_shareBuffer_sbuf_p0_rdat_758,_zz_shareBuffer_sbuf_p0_rdat_759};
  assign _zz_shareBuffer_sbuf_p0_rdat_869 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_870 = {_zz_shareBuffer_sbuf_p0_rdat_871,_zz_shareBuffer_sbuf_p0_rdat_872};
  assign _zz_shareBuffer_sbuf_p0_rdat_984 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_985 = {_zz_shareBuffer_sbuf_p0_rdat_986,_zz_shareBuffer_sbuf_p0_rdat_987};
  assign _zz_shareBuffer_sbuf_p0_rdat_1097 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1098 = {_zz_shareBuffer_sbuf_p0_rdat_1099,_zz_shareBuffer_sbuf_p0_rdat_1100};
  assign _zz_shareBuffer_sbuf_p0_rdat_1211 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1212 = {_zz_shareBuffer_sbuf_p0_rdat_1213,_zz_shareBuffer_sbuf_p0_rdat_1214};
  assign _zz_shareBuffer_sbuf_p0_rdat_1324 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1325 = {_zz_shareBuffer_sbuf_p0_rdat_1326,_zz_shareBuffer_sbuf_p0_rdat_1327};
  assign _zz_shareBuffer_sbuf_p0_rdat_1437 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1438 = {_zz_shareBuffer_sbuf_p0_rdat_1439,_zz_shareBuffer_sbuf_p0_rdat_1440};
  assign _zz_shareBuffer_sbuf_p0_rdat_1549 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1550 = {_zz_shareBuffer_sbuf_p0_rdat_1551,_zz_shareBuffer_sbuf_p0_rdat_1552};
  assign _zz_shareBuffer_sbuf_p0_rdat_1661 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1662 = {_zz_shareBuffer_sbuf_p0_rdat_1663,_zz_shareBuffer_sbuf_p0_rdat_1664};
  assign _zz_shareBuffer_sbuf_p0_rdat_1771 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1772 = {_zz_shareBuffer_sbuf_p0_rdat_1773,_zz_shareBuffer_sbuf_p0_rdat_1774};
  assign _zz_shareBuffer_sbuf_p0_rdat_88 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_89 = {_zz_shareBuffer_sbuf_p0_rdat_90,_zz_shareBuffer_sbuf_p0_rdat_91};
  assign _zz_shareBuffer_sbuf_p0_rdat_197 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_198 = {_zz_shareBuffer_sbuf_p0_rdat_199,_zz_shareBuffer_sbuf_p0_rdat_200};
  assign _zz_shareBuffer_sbuf_p0_rdat_308 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_309 = {_zz_shareBuffer_sbuf_p0_rdat_310,_zz_shareBuffer_sbuf_p0_rdat_311};
  assign _zz_shareBuffer_sbuf_p0_rdat_419 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_420 = {_zz_shareBuffer_sbuf_p0_rdat_421,_zz_shareBuffer_sbuf_p0_rdat_422};
  assign _zz_shareBuffer_sbuf_p0_rdat_532 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_533 = {_zz_shareBuffer_sbuf_p0_rdat_534,_zz_shareBuffer_sbuf_p0_rdat_535};
  assign _zz_shareBuffer_sbuf_p0_rdat_645 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_646 = {_zz_shareBuffer_sbuf_p0_rdat_647,_zz_shareBuffer_sbuf_p0_rdat_648};
  assign _zz_shareBuffer_sbuf_p0_rdat_758 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_759 = {_zz_shareBuffer_sbuf_p0_rdat_760,_zz_shareBuffer_sbuf_p0_rdat_761};
  assign _zz_shareBuffer_sbuf_p0_rdat_871 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_872 = {_zz_shareBuffer_sbuf_p0_rdat_873,_zz_shareBuffer_sbuf_p0_rdat_874};
  assign _zz_shareBuffer_sbuf_p0_rdat_986 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_987 = {_zz_shareBuffer_sbuf_p0_rdat_988,_zz_shareBuffer_sbuf_p0_rdat_989};
  assign _zz_shareBuffer_sbuf_p0_rdat_1099 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1100 = {_zz_shareBuffer_sbuf_p0_rdat_1101,_zz_shareBuffer_sbuf_p0_rdat_1102};
  assign _zz_shareBuffer_sbuf_p0_rdat_1213 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1214 = {_zz_shareBuffer_sbuf_p0_rdat_1215,_zz_shareBuffer_sbuf_p0_rdat_1216};
  assign _zz_shareBuffer_sbuf_p0_rdat_1326 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1327 = {_zz_shareBuffer_sbuf_p0_rdat_1328,_zz_shareBuffer_sbuf_p0_rdat_1329};
  assign _zz_shareBuffer_sbuf_p0_rdat_1439 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1440 = {_zz_shareBuffer_sbuf_p0_rdat_1441,_zz_shareBuffer_sbuf_p0_rdat_1442};
  assign _zz_shareBuffer_sbuf_p0_rdat_1551 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1552 = {_zz_shareBuffer_sbuf_p0_rdat_1553,_zz_shareBuffer_sbuf_p0_rdat_1554};
  assign _zz_shareBuffer_sbuf_p0_rdat_1663 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1664 = {_zz_shareBuffer_sbuf_p0_rdat_1665,_zz_shareBuffer_sbuf_p0_rdat_1666};
  assign _zz_shareBuffer_sbuf_p0_rdat_1773 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1774 = {_zz_shareBuffer_sbuf_p0_rdat_1775,_zz_shareBuffer_sbuf_p0_rdat_1776};
  assign _zz_shareBuffer_sbuf_p0_rdat_90 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_91 = {_zz_shareBuffer_sbuf_p0_rdat_92,_zz_shareBuffer_sbuf_p0_rdat_93};
  assign _zz_shareBuffer_sbuf_p0_rdat_199 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_200 = {_zz_shareBuffer_sbuf_p0_rdat_201,_zz_shareBuffer_sbuf_p0_rdat_202};
  assign _zz_shareBuffer_sbuf_p0_rdat_310 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_311 = {_zz_shareBuffer_sbuf_p0_rdat_312,_zz_shareBuffer_sbuf_p0_rdat_313};
  assign _zz_shareBuffer_sbuf_p0_rdat_421 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_422 = {_zz_shareBuffer_sbuf_p0_rdat_423,_zz_shareBuffer_sbuf_p0_rdat_424};
  assign _zz_shareBuffer_sbuf_p0_rdat_534 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_535 = {_zz_shareBuffer_sbuf_p0_rdat_536,_zz_shareBuffer_sbuf_p0_rdat_537};
  assign _zz_shareBuffer_sbuf_p0_rdat_647 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_648 = {_zz_shareBuffer_sbuf_p0_rdat_649,_zz_shareBuffer_sbuf_p0_rdat_650};
  assign _zz_shareBuffer_sbuf_p0_rdat_760 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_761 = {_zz_shareBuffer_sbuf_p0_rdat_762,_zz_shareBuffer_sbuf_p0_rdat_763};
  assign _zz_shareBuffer_sbuf_p0_rdat_873 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_874 = {_zz_shareBuffer_sbuf_p0_rdat_875,_zz_shareBuffer_sbuf_p0_rdat_876};
  assign _zz_shareBuffer_sbuf_p0_rdat_988 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_989 = {_zz_shareBuffer_sbuf_p0_rdat_990,_zz_shareBuffer_sbuf_p0_rdat_991};
  assign _zz_shareBuffer_sbuf_p0_rdat_1101 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1102 = {_zz_shareBuffer_sbuf_p0_rdat_1103,_zz_shareBuffer_sbuf_p0_rdat_1104};
  assign _zz_shareBuffer_sbuf_p0_rdat_1215 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1216 = {_zz_shareBuffer_sbuf_p0_rdat_1217,_zz_shareBuffer_sbuf_p0_rdat_1218};
  assign _zz_shareBuffer_sbuf_p0_rdat_1328 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1329 = {_zz_shareBuffer_sbuf_p0_rdat_1330,_zz_shareBuffer_sbuf_p0_rdat_1331};
  assign _zz_shareBuffer_sbuf_p0_rdat_1441 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1442 = {_zz_shareBuffer_sbuf_p0_rdat_1443,_zz_shareBuffer_sbuf_p0_rdat_1444};
  assign _zz_shareBuffer_sbuf_p0_rdat_1553 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1554 = {_zz_shareBuffer_sbuf_p0_rdat_1555,_zz_shareBuffer_sbuf_p0_rdat_1556};
  assign _zz_shareBuffer_sbuf_p0_rdat_1665 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1666 = {_zz_shareBuffer_sbuf_p0_rdat_1667,_zz_shareBuffer_sbuf_p0_rdat_1668};
  assign _zz_shareBuffer_sbuf_p0_rdat_1775 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1776 = {_zz_shareBuffer_sbuf_p0_rdat_1777,_zz_shareBuffer_sbuf_p0_rdat_1778};
  assign _zz_shareBuffer_sbuf_p0_rdat_92 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_93 = {_zz_shareBuffer_sbuf_p0_rdat_94,_zz_shareBuffer_sbuf_p0_rdat_95};
  assign _zz_shareBuffer_sbuf_p0_rdat_201 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_202 = {_zz_shareBuffer_sbuf_p0_rdat_203,_zz_shareBuffer_sbuf_p0_rdat_204};
  assign _zz_shareBuffer_sbuf_p0_rdat_312 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_313 = {_zz_shareBuffer_sbuf_p0_rdat_314,_zz_shareBuffer_sbuf_p0_rdat_315};
  assign _zz_shareBuffer_sbuf_p0_rdat_423 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_424 = {_zz_shareBuffer_sbuf_p0_rdat_425,_zz_shareBuffer_sbuf_p0_rdat_426};
  assign _zz_shareBuffer_sbuf_p0_rdat_536 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_537 = {_zz_shareBuffer_sbuf_p0_rdat_538,_zz_shareBuffer_sbuf_p0_rdat_539};
  assign _zz_shareBuffer_sbuf_p0_rdat_649 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_650 = {_zz_shareBuffer_sbuf_p0_rdat_651,_zz_shareBuffer_sbuf_p0_rdat_652};
  assign _zz_shareBuffer_sbuf_p0_rdat_762 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_763 = {_zz_shareBuffer_sbuf_p0_rdat_764,_zz_shareBuffer_sbuf_p0_rdat_765};
  assign _zz_shareBuffer_sbuf_p0_rdat_875 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_876 = {_zz_shareBuffer_sbuf_p0_rdat_877,_zz_shareBuffer_sbuf_p0_rdat_878};
  assign _zz_shareBuffer_sbuf_p0_rdat_990 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_991 = {_zz_shareBuffer_sbuf_p0_rdat_992,_zz_shareBuffer_sbuf_p0_rdat_993};
  assign _zz_shareBuffer_sbuf_p0_rdat_1103 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1104 = {_zz_shareBuffer_sbuf_p0_rdat_1105,_zz_shareBuffer_sbuf_p0_rdat_1106};
  assign _zz_shareBuffer_sbuf_p0_rdat_1217 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1218 = {_zz_shareBuffer_sbuf_p0_rdat_1219,_zz_shareBuffer_sbuf_p0_rdat_1220};
  assign _zz_shareBuffer_sbuf_p0_rdat_1330 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1331 = {_zz_shareBuffer_sbuf_p0_rdat_1332,_zz_shareBuffer_sbuf_p0_rdat_1333};
  assign _zz_shareBuffer_sbuf_p0_rdat_1443 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1444 = {_zz_shareBuffer_sbuf_p0_rdat_1445,_zz_shareBuffer_sbuf_p0_rdat_1446};
  assign _zz_shareBuffer_sbuf_p0_rdat_1555 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1556 = {_zz_shareBuffer_sbuf_p0_rdat_1557,_zz_shareBuffer_sbuf_p0_rdat_1558};
  assign _zz_shareBuffer_sbuf_p0_rdat_1667 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1668 = {_zz_shareBuffer_sbuf_p0_rdat_1669,_zz_shareBuffer_sbuf_p0_rdat_1670};
  assign _zz_shareBuffer_sbuf_p0_rdat_1777 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1778 = {_zz_shareBuffer_sbuf_p0_rdat_1779,_zz_shareBuffer_sbuf_p0_rdat_1780};
  assign _zz_shareBuffer_sbuf_p0_rdat_94 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_95 = {_zz_shareBuffer_sbuf_p0_rdat_96,_zz_shareBuffer_sbuf_p0_rdat_97};
  assign _zz_shareBuffer_sbuf_p0_rdat_203 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_204 = {_zz_shareBuffer_sbuf_p0_rdat_205,_zz_shareBuffer_sbuf_p0_rdat_206};
  assign _zz_shareBuffer_sbuf_p0_rdat_314 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_315 = {_zz_shareBuffer_sbuf_p0_rdat_316,_zz_shareBuffer_sbuf_p0_rdat_317};
  assign _zz_shareBuffer_sbuf_p0_rdat_425 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_426 = {_zz_shareBuffer_sbuf_p0_rdat_427,_zz_shareBuffer_sbuf_p0_rdat_428};
  assign _zz_shareBuffer_sbuf_p0_rdat_538 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_539 = {_zz_shareBuffer_sbuf_p0_rdat_540,_zz_shareBuffer_sbuf_p0_rdat_541};
  assign _zz_shareBuffer_sbuf_p0_rdat_651 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_652 = {_zz_shareBuffer_sbuf_p0_rdat_653,_zz_shareBuffer_sbuf_p0_rdat_654};
  assign _zz_shareBuffer_sbuf_p0_rdat_764 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_765 = {_zz_shareBuffer_sbuf_p0_rdat_766,_zz_shareBuffer_sbuf_p0_rdat_767};
  assign _zz_shareBuffer_sbuf_p0_rdat_877 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_878 = {_zz_shareBuffer_sbuf_p0_rdat_879,_zz_shareBuffer_sbuf_p0_rdat_880};
  assign _zz_shareBuffer_sbuf_p0_rdat_992 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_993 = {_zz_shareBuffer_sbuf_p0_rdat_994,_zz_shareBuffer_sbuf_p0_rdat_995};
  assign _zz_shareBuffer_sbuf_p0_rdat_1105 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1106 = {_zz_shareBuffer_sbuf_p0_rdat_1107,_zz_shareBuffer_sbuf_p0_rdat_1108};
  assign _zz_shareBuffer_sbuf_p0_rdat_1219 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1220 = {_zz_shareBuffer_sbuf_p0_rdat_1221,_zz_shareBuffer_sbuf_p0_rdat_1222};
  assign _zz_shareBuffer_sbuf_p0_rdat_1332 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1333 = {_zz_shareBuffer_sbuf_p0_rdat_1334,_zz_shareBuffer_sbuf_p0_rdat_1335};
  assign _zz_shareBuffer_sbuf_p0_rdat_1445 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1446 = {_zz_shareBuffer_sbuf_p0_rdat_1447,_zz_shareBuffer_sbuf_p0_rdat_1448};
  assign _zz_shareBuffer_sbuf_p0_rdat_1557 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1558 = {_zz_shareBuffer_sbuf_p0_rdat_1559,_zz_shareBuffer_sbuf_p0_rdat_1560};
  assign _zz_shareBuffer_sbuf_p0_rdat_1669 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1670 = {_zz_shareBuffer_sbuf_p0_rdat_1671,_zz_shareBuffer_sbuf_p0_rdat_1672};
  assign _zz_shareBuffer_sbuf_p0_rdat_1779 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1780 = {_zz_shareBuffer_sbuf_p0_rdat_1781,_zz_shareBuffer_sbuf_p0_rdat_1782};
  assign _zz_shareBuffer_sbuf_p0_rdat_96 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_97 = {_zz_shareBuffer_sbuf_p0_rdat_98,_zz_shareBuffer_sbuf_p0_rdat_99};
  assign _zz_shareBuffer_sbuf_p0_rdat_205 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_206 = {_zz_shareBuffer_sbuf_p0_rdat_207,_zz_shareBuffer_sbuf_p0_rdat_208};
  assign _zz_shareBuffer_sbuf_p0_rdat_316 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_317 = {_zz_shareBuffer_sbuf_p0_rdat_318,_zz_shareBuffer_sbuf_p0_rdat_319};
  assign _zz_shareBuffer_sbuf_p0_rdat_427 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_428 = {_zz_shareBuffer_sbuf_p0_rdat_429,_zz_shareBuffer_sbuf_p0_rdat_430};
  assign _zz_shareBuffer_sbuf_p0_rdat_540 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_541 = {_zz_shareBuffer_sbuf_p0_rdat_542,_zz_shareBuffer_sbuf_p0_rdat_543};
  assign _zz_shareBuffer_sbuf_p0_rdat_653 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_654 = {_zz_shareBuffer_sbuf_p0_rdat_655,_zz_shareBuffer_sbuf_p0_rdat_656};
  assign _zz_shareBuffer_sbuf_p0_rdat_766 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_767 = {_zz_shareBuffer_sbuf_p0_rdat_768,_zz_shareBuffer_sbuf_p0_rdat_769};
  assign _zz_shareBuffer_sbuf_p0_rdat_879 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_880 = {_zz_shareBuffer_sbuf_p0_rdat_881,_zz_shareBuffer_sbuf_p0_rdat_882};
  assign _zz_shareBuffer_sbuf_p0_rdat_994 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_995 = {_zz_shareBuffer_sbuf_p0_rdat_996,_zz_shareBuffer_sbuf_p0_rdat_997};
  assign _zz_shareBuffer_sbuf_p0_rdat_1107 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1108 = {_zz_shareBuffer_sbuf_p0_rdat_1109,_zz_shareBuffer_sbuf_p0_rdat_1110};
  assign _zz_shareBuffer_sbuf_p0_rdat_1221 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1222 = {_zz_shareBuffer_sbuf_p0_rdat_1223,_zz_shareBuffer_sbuf_p0_rdat_1224};
  assign _zz_shareBuffer_sbuf_p0_rdat_1334 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1335 = {_zz_shareBuffer_sbuf_p0_rdat_1336,_zz_shareBuffer_sbuf_p0_rdat_1337};
  assign _zz_shareBuffer_sbuf_p0_rdat_1447 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1448 = {_zz_shareBuffer_sbuf_p0_rdat_1449,_zz_shareBuffer_sbuf_p0_rdat_1450};
  assign _zz_shareBuffer_sbuf_p0_rdat_1559 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1560 = {_zz_shareBuffer_sbuf_p0_rdat_1561,_zz_shareBuffer_sbuf_p0_rdat_1562};
  assign _zz_shareBuffer_sbuf_p0_rdat_1671 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1672 = {_zz_shareBuffer_sbuf_p0_rdat_1673,_zz_shareBuffer_sbuf_p0_rdat_1674};
  assign _zz_shareBuffer_sbuf_p0_rdat_1781 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1782 = {_zz_shareBuffer_sbuf_p0_rdat_1783,_zz_shareBuffer_sbuf_p0_rdat_1784};
  assign _zz_shareBuffer_sbuf_p0_rdat_98 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_99 = {_zz_shareBuffer_sbuf_p0_rdat_100,_zz_shareBuffer_sbuf_p0_rdat_101};
  assign _zz_shareBuffer_sbuf_p0_rdat_207 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_208 = {_zz_shareBuffer_sbuf_p0_rdat_209,_zz_shareBuffer_sbuf_p0_rdat_210};
  assign _zz_shareBuffer_sbuf_p0_rdat_318 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_319 = {_zz_shareBuffer_sbuf_p0_rdat_320,_zz_shareBuffer_sbuf_p0_rdat_321};
  assign _zz_shareBuffer_sbuf_p0_rdat_429 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_430 = {_zz_shareBuffer_sbuf_p0_rdat_431,_zz_shareBuffer_sbuf_p0_rdat_432};
  assign _zz_shareBuffer_sbuf_p0_rdat_542 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_543 = {_zz_shareBuffer_sbuf_p0_rdat_544,_zz_shareBuffer_sbuf_p0_rdat_545};
  assign _zz_shareBuffer_sbuf_p0_rdat_655 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_656 = {_zz_shareBuffer_sbuf_p0_rdat_657,_zz_shareBuffer_sbuf_p0_rdat_658};
  assign _zz_shareBuffer_sbuf_p0_rdat_768 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_769 = {_zz_shareBuffer_sbuf_p0_rdat_770,_zz_shareBuffer_sbuf_p0_rdat_771};
  assign _zz_shareBuffer_sbuf_p0_rdat_881 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_882 = {_zz_shareBuffer_sbuf_p0_rdat_883,_zz_shareBuffer_sbuf_p0_rdat_884};
  assign _zz_shareBuffer_sbuf_p0_rdat_996 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_997 = {_zz_shareBuffer_sbuf_p0_rdat_998,_zz_shareBuffer_sbuf_p0_rdat_999};
  assign _zz_shareBuffer_sbuf_p0_rdat_1109 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1110 = {_zz_shareBuffer_sbuf_p0_rdat_1111,_zz_shareBuffer_sbuf_p0_rdat_1112};
  assign _zz_shareBuffer_sbuf_p0_rdat_1223 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1224 = {_zz_shareBuffer_sbuf_p0_rdat_1225,_zz_shareBuffer_sbuf_p0_rdat_1226};
  assign _zz_shareBuffer_sbuf_p0_rdat_1336 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1337 = {_zz_shareBuffer_sbuf_p0_rdat_1338,_zz_shareBuffer_sbuf_p0_rdat_1339};
  assign _zz_shareBuffer_sbuf_p0_rdat_1449 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1450 = {_zz_shareBuffer_sbuf_p0_rdat_1451,_zz_shareBuffer_sbuf_p0_rdat_1452};
  assign _zz_shareBuffer_sbuf_p0_rdat_1561 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1562 = {_zz_shareBuffer_sbuf_p0_rdat_1563,_zz_shareBuffer_sbuf_p0_rdat_1564};
  assign _zz_shareBuffer_sbuf_p0_rdat_1673 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1674 = {_zz_shareBuffer_sbuf_p0_rdat_1675,_zz_shareBuffer_sbuf_p0_rdat_1676};
  assign _zz_shareBuffer_sbuf_p0_rdat_1783 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1784 = {_zz_shareBuffer_sbuf_p0_rdat_1785,_zz_shareBuffer_sbuf_p0_rdat_1786};
  assign _zz_shareBuffer_sbuf_p0_rdat_100 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_101 = {_zz_shareBuffer_sbuf_p0_rdat_102,_zz_shareBuffer_sbuf_p0_rdat_103};
  assign _zz_shareBuffer_sbuf_p0_rdat_209 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_210 = {_zz_shareBuffer_sbuf_p0_rdat_211,_zz_shareBuffer_sbuf_p0_rdat_212};
  assign _zz_shareBuffer_sbuf_p0_rdat_320 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_321 = {_zz_shareBuffer_sbuf_p0_rdat_322,_zz_shareBuffer_sbuf_p0_rdat_323};
  assign _zz_shareBuffer_sbuf_p0_rdat_431 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_432 = {_zz_shareBuffer_sbuf_p0_rdat_433,_zz_shareBuffer_sbuf_p0_rdat_434};
  assign _zz_shareBuffer_sbuf_p0_rdat_544 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_545 = {_zz_shareBuffer_sbuf_p0_rdat_546,_zz_shareBuffer_sbuf_p0_rdat_547};
  assign _zz_shareBuffer_sbuf_p0_rdat_657 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_658 = {_zz_shareBuffer_sbuf_p0_rdat_659,_zz_shareBuffer_sbuf_p0_rdat_660};
  assign _zz_shareBuffer_sbuf_p0_rdat_770 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_771 = {_zz_shareBuffer_sbuf_p0_rdat_772,_zz_shareBuffer_sbuf_p0_rdat_773};
  assign _zz_shareBuffer_sbuf_p0_rdat_883 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_884 = {_zz_shareBuffer_sbuf_p0_rdat_885,_zz_shareBuffer_sbuf_p0_rdat_886};
  assign _zz_shareBuffer_sbuf_p0_rdat_998 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_999 = {_zz_shareBuffer_sbuf_p0_rdat_1000,_zz_shareBuffer_sbuf_p0_rdat_1001};
  assign _zz_shareBuffer_sbuf_p0_rdat_1111 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1112 = {_zz_shareBuffer_sbuf_p0_rdat_1113,_zz_shareBuffer_sbuf_p0_rdat_1114};
  assign _zz_shareBuffer_sbuf_p0_rdat_1225 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1226 = {_zz_shareBuffer_sbuf_p0_rdat_1227,_zz_shareBuffer_sbuf_p0_rdat_1228};
  assign _zz_shareBuffer_sbuf_p0_rdat_1338 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1339 = {_zz_shareBuffer_sbuf_p0_rdat_1340,_zz_shareBuffer_sbuf_p0_rdat_1341};
  assign _zz_shareBuffer_sbuf_p0_rdat_1451 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1452 = {_zz_shareBuffer_sbuf_p0_rdat_1453,_zz_shareBuffer_sbuf_p0_rdat_1454};
  assign _zz_shareBuffer_sbuf_p0_rdat_1563 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1564 = {_zz_shareBuffer_sbuf_p0_rdat_1565,_zz_shareBuffer_sbuf_p0_rdat_1566};
  assign _zz_shareBuffer_sbuf_p0_rdat_1675 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1676 = {_zz_shareBuffer_sbuf_p0_rdat_1677,_zz_shareBuffer_sbuf_p0_rdat_1678};
  assign _zz_shareBuffer_sbuf_p0_rdat_1785 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1786 = {_zz_shareBuffer_sbuf_p0_rdat_1787,_zz_shareBuffer_sbuf_p0_rdat_1788};
  assign _zz_shareBuffer_sbuf_p0_rdat_102 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_103 = {shareBuffer_sbuf_p0_re_norm_d1_0,{_zz_shareBuffer_sbuf_p0_rdat_104,_zz_shareBuffer_sbuf_p0_rdat_105}};
  assign _zz_shareBuffer_sbuf_p0_rdat_211 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_212 = {shareBuffer_sbuf_p0_re_norm_d1_1,{_zz_shareBuffer_sbuf_p0_rdat_213,_zz_shareBuffer_sbuf_p0_rdat_214}};
  assign _zz_shareBuffer_sbuf_p0_rdat_322 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_323 = {shareBuffer_sbuf_p0_re_norm_d1_2,{_zz_shareBuffer_sbuf_p0_rdat_324,_zz_shareBuffer_sbuf_p0_rdat_325}};
  assign _zz_shareBuffer_sbuf_p0_rdat_433 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_434 = {shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_435,_zz_shareBuffer_sbuf_p0_rdat_436}};
  assign _zz_shareBuffer_sbuf_p0_rdat_546 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_547 = {shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_548,_zz_shareBuffer_sbuf_p0_rdat_549}};
  assign _zz_shareBuffer_sbuf_p0_rdat_659 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_660 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_661,_zz_shareBuffer_sbuf_p0_rdat_662}};
  assign _zz_shareBuffer_sbuf_p0_rdat_772 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_773 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_774,_zz_shareBuffer_sbuf_p0_rdat_775}};
  assign _zz_shareBuffer_sbuf_p0_rdat_885 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_886 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_887,_zz_shareBuffer_sbuf_p0_rdat_888}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1000 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_1001 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_1002,_zz_shareBuffer_sbuf_p0_rdat_1003}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1113 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1114 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1115,_zz_shareBuffer_sbuf_p0_rdat_1116}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1227 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1228 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1229,_zz_shareBuffer_sbuf_p0_rdat_1230}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1340 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1341 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1342,_zz_shareBuffer_sbuf_p0_rdat_1343}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1453 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1454 = {shareBuffer_sbuf_p0_re_norm_d1_12,{_zz_shareBuffer_sbuf_p0_rdat_1455,_zz_shareBuffer_sbuf_p0_rdat_1456}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1565 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1566 = {shareBuffer_sbuf_p0_re_norm_d1_13,{_zz_shareBuffer_sbuf_p0_rdat_1567,_zz_shareBuffer_sbuf_p0_rdat_1568}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1677 = shareBuffer_sbuf_p0_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p0_rdat_1678 = {shareBuffer_sbuf_p0_re_norm_d1_14,shareBuffer_sbuf_p0_re_norm_d1_14};
  assign _zz_shareBuffer_sbuf_p0_rdat_1787 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_1788 = shareBuffer_sbuf_p0_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p0_rdat_104 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_105 = {shareBuffer_sbuf_p0_re_norm_d1_0,{_zz_shareBuffer_sbuf_p0_rdat_106,_zz_shareBuffer_sbuf_p0_rdat_107}};
  assign _zz_shareBuffer_sbuf_p0_rdat_213 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_214 = {shareBuffer_sbuf_p0_re_norm_d1_1,{_zz_shareBuffer_sbuf_p0_rdat_215,_zz_shareBuffer_sbuf_p0_rdat_216}};
  assign _zz_shareBuffer_sbuf_p0_rdat_324 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_325 = {shareBuffer_sbuf_p0_re_norm_d1_2,{_zz_shareBuffer_sbuf_p0_rdat_326,_zz_shareBuffer_sbuf_p0_rdat_327}};
  assign _zz_shareBuffer_sbuf_p0_rdat_435 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_436 = {shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_437,_zz_shareBuffer_sbuf_p0_rdat_438}};
  assign _zz_shareBuffer_sbuf_p0_rdat_548 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_549 = {shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_550,_zz_shareBuffer_sbuf_p0_rdat_551}};
  assign _zz_shareBuffer_sbuf_p0_rdat_661 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_662 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_663,_zz_shareBuffer_sbuf_p0_rdat_664}};
  assign _zz_shareBuffer_sbuf_p0_rdat_774 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_775 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_776,_zz_shareBuffer_sbuf_p0_rdat_777}};
  assign _zz_shareBuffer_sbuf_p0_rdat_887 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_888 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_889,_zz_shareBuffer_sbuf_p0_rdat_890}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1002 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_1003 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_1004,_zz_shareBuffer_sbuf_p0_rdat_1005}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1115 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1116 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1117,_zz_shareBuffer_sbuf_p0_rdat_1118}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1229 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1230 = {shareBuffer_sbuf_p0_re_norm_d1_10,{_zz_shareBuffer_sbuf_p0_rdat_1231,_zz_shareBuffer_sbuf_p0_rdat_1232}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1342 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1343 = {shareBuffer_sbuf_p0_re_norm_d1_11,{_zz_shareBuffer_sbuf_p0_rdat_1344,_zz_shareBuffer_sbuf_p0_rdat_1345}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1455 = shareBuffer_sbuf_p0_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p0_rdat_1456 = {shareBuffer_sbuf_p0_re_norm_d1_12,shareBuffer_sbuf_p0_re_norm_d1_12};
  assign _zz_shareBuffer_sbuf_p0_rdat_1567 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_1568 = shareBuffer_sbuf_p0_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p0_rdat_106 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_107 = {shareBuffer_sbuf_p0_re_norm_d1_0,{_zz_shareBuffer_sbuf_p0_rdat_108,_zz_shareBuffer_sbuf_p0_rdat_109}};
  assign _zz_shareBuffer_sbuf_p0_rdat_215 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_216 = {shareBuffer_sbuf_p0_re_norm_d1_1,{_zz_shareBuffer_sbuf_p0_rdat_217,_zz_shareBuffer_sbuf_p0_rdat_218}};
  assign _zz_shareBuffer_sbuf_p0_rdat_326 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_327 = {shareBuffer_sbuf_p0_re_norm_d1_2,{_zz_shareBuffer_sbuf_p0_rdat_328,_zz_shareBuffer_sbuf_p0_rdat_329}};
  assign _zz_shareBuffer_sbuf_p0_rdat_437 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_438 = {shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_439,_zz_shareBuffer_sbuf_p0_rdat_440}};
  assign _zz_shareBuffer_sbuf_p0_rdat_550 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_551 = {shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_552,_zz_shareBuffer_sbuf_p0_rdat_553}};
  assign _zz_shareBuffer_sbuf_p0_rdat_663 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_664 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_665,_zz_shareBuffer_sbuf_p0_rdat_666}};
  assign _zz_shareBuffer_sbuf_p0_rdat_776 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_777 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_778,_zz_shareBuffer_sbuf_p0_rdat_779}};
  assign _zz_shareBuffer_sbuf_p0_rdat_889 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_890 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_891,_zz_shareBuffer_sbuf_p0_rdat_892}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1004 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_1005 = {shareBuffer_sbuf_p0_re_norm_d1_8,{_zz_shareBuffer_sbuf_p0_rdat_1006,_zz_shareBuffer_sbuf_p0_rdat_1007}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1117 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1118 = {shareBuffer_sbuf_p0_re_norm_d1_9,{_zz_shareBuffer_sbuf_p0_rdat_1119,_zz_shareBuffer_sbuf_p0_rdat_1120}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1231 = shareBuffer_sbuf_p0_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p0_rdat_1232 = {shareBuffer_sbuf_p0_re_norm_d1_10,shareBuffer_sbuf_p0_re_norm_d1_10};
  assign _zz_shareBuffer_sbuf_p0_rdat_1344 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_1345 = shareBuffer_sbuf_p0_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p0_rdat_108 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_109 = {shareBuffer_sbuf_p0_re_norm_d1_0,{_zz_shareBuffer_sbuf_p0_rdat_110,_zz_shareBuffer_sbuf_p0_rdat_111}};
  assign _zz_shareBuffer_sbuf_p0_rdat_217 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_218 = {shareBuffer_sbuf_p0_re_norm_d1_1,{_zz_shareBuffer_sbuf_p0_rdat_219,_zz_shareBuffer_sbuf_p0_rdat_220}};
  assign _zz_shareBuffer_sbuf_p0_rdat_328 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_329 = {shareBuffer_sbuf_p0_re_norm_d1_2,{_zz_shareBuffer_sbuf_p0_rdat_330,_zz_shareBuffer_sbuf_p0_rdat_331}};
  assign _zz_shareBuffer_sbuf_p0_rdat_439 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_440 = {shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_441,_zz_shareBuffer_sbuf_p0_rdat_442}};
  assign _zz_shareBuffer_sbuf_p0_rdat_552 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_553 = {shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_554,_zz_shareBuffer_sbuf_p0_rdat_555}};
  assign _zz_shareBuffer_sbuf_p0_rdat_665 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_666 = {shareBuffer_sbuf_p0_re_norm_d1_5,{_zz_shareBuffer_sbuf_p0_rdat_667,_zz_shareBuffer_sbuf_p0_rdat_668}};
  assign _zz_shareBuffer_sbuf_p0_rdat_778 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_779 = {shareBuffer_sbuf_p0_re_norm_d1_6,{_zz_shareBuffer_sbuf_p0_rdat_780,_zz_shareBuffer_sbuf_p0_rdat_781}};
  assign _zz_shareBuffer_sbuf_p0_rdat_891 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_892 = {shareBuffer_sbuf_p0_re_norm_d1_7,{_zz_shareBuffer_sbuf_p0_rdat_893,_zz_shareBuffer_sbuf_p0_rdat_894}};
  assign _zz_shareBuffer_sbuf_p0_rdat_1006 = shareBuffer_sbuf_p0_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p0_rdat_1007 = {shareBuffer_sbuf_p0_re_norm_d1_8,shareBuffer_sbuf_p0_re_norm_d1_8};
  assign _zz_shareBuffer_sbuf_p0_rdat_1119 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_1120 = shareBuffer_sbuf_p0_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p0_rdat_110 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_111 = {shareBuffer_sbuf_p0_re_norm_d1_0,{shareBuffer_sbuf_p0_re_norm_d1_0,{_zz_shareBuffer_sbuf_p0_rdat_112,_zz_shareBuffer_sbuf_p0_rdat_113}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_219 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_220 = {shareBuffer_sbuf_p0_re_norm_d1_1,{shareBuffer_sbuf_p0_re_norm_d1_1,{_zz_shareBuffer_sbuf_p0_rdat_221,_zz_shareBuffer_sbuf_p0_rdat_222}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_330 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_331 = {shareBuffer_sbuf_p0_re_norm_d1_2,{shareBuffer_sbuf_p0_re_norm_d1_2,{_zz_shareBuffer_sbuf_p0_rdat_332,_zz_shareBuffer_sbuf_p0_rdat_333}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_441 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_442 = {shareBuffer_sbuf_p0_re_norm_d1_3,{shareBuffer_sbuf_p0_re_norm_d1_3,{_zz_shareBuffer_sbuf_p0_rdat_443,_zz_shareBuffer_sbuf_p0_rdat_444}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_554 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_555 = {shareBuffer_sbuf_p0_re_norm_d1_4,{shareBuffer_sbuf_p0_re_norm_d1_4,{_zz_shareBuffer_sbuf_p0_rdat_556,_zz_shareBuffer_sbuf_p0_rdat_557}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_667 = shareBuffer_sbuf_p0_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p0_rdat_668 = {shareBuffer_sbuf_p0_re_norm_d1_5,{shareBuffer_sbuf_p0_re_norm_d1_5,shareBuffer_sbuf_p0_re_norm_d1_5}};
  assign _zz_shareBuffer_sbuf_p0_rdat_780 = shareBuffer_sbuf_p0_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p0_rdat_781 = {shareBuffer_sbuf_p0_re_norm_d1_6,shareBuffer_sbuf_p0_re_norm_d1_6};
  assign _zz_shareBuffer_sbuf_p0_rdat_893 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_894 = shareBuffer_sbuf_p0_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p0_rdat_112 = shareBuffer_sbuf_p0_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p0_rdat_113 = {shareBuffer_sbuf_p0_re_norm_d1_0,{shareBuffer_sbuf_p0_re_norm_d1_0,{shareBuffer_sbuf_p0_re_norm_d1_0,shareBuffer_sbuf_p0_re_norm_d1_0}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_221 = shareBuffer_sbuf_p0_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p0_rdat_222 = {shareBuffer_sbuf_p0_re_norm_d1_1,{shareBuffer_sbuf_p0_re_norm_d1_1,{shareBuffer_sbuf_p0_re_norm_d1_1,shareBuffer_sbuf_p0_re_norm_d1_1}}};
  assign _zz_shareBuffer_sbuf_p0_rdat_332 = shareBuffer_sbuf_p0_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p0_rdat_333 = {shareBuffer_sbuf_p0_re_norm_d1_2,{shareBuffer_sbuf_p0_re_norm_d1_2,shareBuffer_sbuf_p0_re_norm_d1_2}};
  assign _zz_shareBuffer_sbuf_p0_rdat_443 = shareBuffer_sbuf_p0_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p0_rdat_444 = {shareBuffer_sbuf_p0_re_norm_d1_3,shareBuffer_sbuf_p0_re_norm_d1_3};
  assign _zz_shareBuffer_sbuf_p0_rdat_556 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p0_rdat_557 = shareBuffer_sbuf_p0_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat = (((_zz_shareBuffer_sbuf_p1_rdat_1 | _zz_shareBuffer_sbuf_p1_rdat_895) | (_zz_shareBuffer_sbuf_p1_rdat_1008 & shareBuffer_sbuf_rdat_9)) | ({_zz_shareBuffer_sbuf_p1_rdat_1121,_zz_shareBuffer_sbuf_p1_rdat_1122} & shareBuffer_sbuf_rdat_10));
  assign _zz_shareBuffer_sbuf_p1_rdat_1233 = ({shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1234,_zz_shareBuffer_sbuf_p1_rdat_1235}} & shareBuffer_sbuf_rdat_11);
  assign _zz_shareBuffer_sbuf_p1_rdat_1346 = {shareBuffer_sbuf_p1_re_norm_d1_12,{shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1347,_zz_shareBuffer_sbuf_p1_rdat_1348}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1457 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1458 = {shareBuffer_sbuf_p1_re_norm_d1_13,{shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1459,_zz_shareBuffer_sbuf_p1_rdat_1460}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1569 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1570 = {shareBuffer_sbuf_p1_re_norm_d1_14,{shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1571,_zz_shareBuffer_sbuf_p1_rdat_1572}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1679 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1680 = {shareBuffer_sbuf_p1_re_norm_d1_15,{shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1681,_zz_shareBuffer_sbuf_p1_rdat_1682}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1 = ((_zz_shareBuffer_sbuf_p1_rdat_2 | _zz_shareBuffer_sbuf_p1_rdat_669) | (_zz_shareBuffer_sbuf_p1_rdat_782 & shareBuffer_sbuf_rdat_7));
  assign _zz_shareBuffer_sbuf_p1_rdat_895 = ({_zz_shareBuffer_sbuf_p1_rdat_896,_zz_shareBuffer_sbuf_p1_rdat_897} & shareBuffer_sbuf_rdat_8);
  assign _zz_shareBuffer_sbuf_p1_rdat_1008 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1009,_zz_shareBuffer_sbuf_p1_rdat_1010}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1121 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1122 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1123,_zz_shareBuffer_sbuf_p1_rdat_1124}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1234 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1235 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1236,_zz_shareBuffer_sbuf_p1_rdat_1237}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1347 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1348 = {shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1349,_zz_shareBuffer_sbuf_p1_rdat_1350}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1459 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1460 = {shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1461,_zz_shareBuffer_sbuf_p1_rdat_1462}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1571 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1572 = {shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1573,_zz_shareBuffer_sbuf_p1_rdat_1574}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1681 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1682 = {shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1683,_zz_shareBuffer_sbuf_p1_rdat_1684}};
  assign _zz_shareBuffer_sbuf_p1_rdat_2 = ((_zz_shareBuffer_sbuf_p1_rdat_3 | _zz_shareBuffer_sbuf_p1_rdat_445) | (_zz_shareBuffer_sbuf_p1_rdat_558 & shareBuffer_sbuf_rdat_5));
  assign _zz_shareBuffer_sbuf_p1_rdat_669 = ({_zz_shareBuffer_sbuf_p1_rdat_670,_zz_shareBuffer_sbuf_p1_rdat_671} & shareBuffer_sbuf_rdat_6);
  assign _zz_shareBuffer_sbuf_p1_rdat_782 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_783,_zz_shareBuffer_sbuf_p1_rdat_784}};
  assign _zz_shareBuffer_sbuf_p1_rdat_896 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_897 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_898,_zz_shareBuffer_sbuf_p1_rdat_899}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1009 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1010 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1011,_zz_shareBuffer_sbuf_p1_rdat_1012}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1123 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1124 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1125,_zz_shareBuffer_sbuf_p1_rdat_1126}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1236 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1237 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1238,_zz_shareBuffer_sbuf_p1_rdat_1239}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1349 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1350 = {shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1351,_zz_shareBuffer_sbuf_p1_rdat_1352}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1461 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1462 = {shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1463,_zz_shareBuffer_sbuf_p1_rdat_1464}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1573 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1574 = {shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1575,_zz_shareBuffer_sbuf_p1_rdat_1576}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1683 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1684 = {shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1685,_zz_shareBuffer_sbuf_p1_rdat_1686}};
  assign _zz_shareBuffer_sbuf_p1_rdat_3 = ((_zz_shareBuffer_sbuf_p1_rdat_4 | _zz_shareBuffer_sbuf_p1_rdat_223) | (_zz_shareBuffer_sbuf_p1_rdat_334 & shareBuffer_sbuf_rdat_3));
  assign _zz_shareBuffer_sbuf_p1_rdat_445 = ({_zz_shareBuffer_sbuf_p1_rdat_446,_zz_shareBuffer_sbuf_p1_rdat_447} & shareBuffer_sbuf_rdat_4);
  assign _zz_shareBuffer_sbuf_p1_rdat_558 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_559,_zz_shareBuffer_sbuf_p1_rdat_560}};
  assign _zz_shareBuffer_sbuf_p1_rdat_670 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_671 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_672,_zz_shareBuffer_sbuf_p1_rdat_673}};
  assign _zz_shareBuffer_sbuf_p1_rdat_783 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_784 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_785,_zz_shareBuffer_sbuf_p1_rdat_786}};
  assign _zz_shareBuffer_sbuf_p1_rdat_898 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_899 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_900,_zz_shareBuffer_sbuf_p1_rdat_901}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1011 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1012 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1013,_zz_shareBuffer_sbuf_p1_rdat_1014}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1125 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1126 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1127,_zz_shareBuffer_sbuf_p1_rdat_1128}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1238 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1239 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1240,_zz_shareBuffer_sbuf_p1_rdat_1241}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1351 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1352 = {shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1353,_zz_shareBuffer_sbuf_p1_rdat_1354}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1463 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1464 = {shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1465,_zz_shareBuffer_sbuf_p1_rdat_1466}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1575 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1576 = {shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1577,_zz_shareBuffer_sbuf_p1_rdat_1578}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1685 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1686 = {shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1687,_zz_shareBuffer_sbuf_p1_rdat_1688}};
  assign _zz_shareBuffer_sbuf_p1_rdat_4 = ((_zz_shareBuffer_sbuf_p1_rdat_5 & shareBuffer_sbuf_rdat_0) | (_zz_shareBuffer_sbuf_p1_rdat_114 & shareBuffer_sbuf_rdat_1));
  assign _zz_shareBuffer_sbuf_p1_rdat_223 = ({_zz_shareBuffer_sbuf_p1_rdat_224,_zz_shareBuffer_sbuf_p1_rdat_225} & shareBuffer_sbuf_rdat_2);
  assign _zz_shareBuffer_sbuf_p1_rdat_334 = {shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_335,_zz_shareBuffer_sbuf_p1_rdat_336}};
  assign _zz_shareBuffer_sbuf_p1_rdat_446 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_447 = {shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_448,_zz_shareBuffer_sbuf_p1_rdat_449}};
  assign _zz_shareBuffer_sbuf_p1_rdat_559 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_560 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_561,_zz_shareBuffer_sbuf_p1_rdat_562}};
  assign _zz_shareBuffer_sbuf_p1_rdat_672 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_673 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_674,_zz_shareBuffer_sbuf_p1_rdat_675}};
  assign _zz_shareBuffer_sbuf_p1_rdat_785 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_786 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_787,_zz_shareBuffer_sbuf_p1_rdat_788}};
  assign _zz_shareBuffer_sbuf_p1_rdat_900 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_901 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_902,_zz_shareBuffer_sbuf_p1_rdat_903}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1013 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1014 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1015,_zz_shareBuffer_sbuf_p1_rdat_1016}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1127 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1128 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1129,_zz_shareBuffer_sbuf_p1_rdat_1130}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1240 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1241 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1242,_zz_shareBuffer_sbuf_p1_rdat_1243}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1353 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1354 = {shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1355,_zz_shareBuffer_sbuf_p1_rdat_1356}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1465 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1466 = {shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1467,_zz_shareBuffer_sbuf_p1_rdat_1468}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1577 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1578 = {shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1579,_zz_shareBuffer_sbuf_p1_rdat_1580}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1687 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1688 = {shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1689,_zz_shareBuffer_sbuf_p1_rdat_1690}};
  assign _zz_shareBuffer_sbuf_p1_rdat_5 = {_zz_shareBuffer_sbuf_p1_rdat_6,_zz_shareBuffer_sbuf_p1_rdat_7};
  assign _zz_shareBuffer_sbuf_p1_rdat_114 = {_zz_shareBuffer_sbuf_p1_rdat_115,_zz_shareBuffer_sbuf_p1_rdat_116};
  assign _zz_shareBuffer_sbuf_p1_rdat_224 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_225 = {_zz_shareBuffer_sbuf_p1_rdat_226,_zz_shareBuffer_sbuf_p1_rdat_227};
  assign _zz_shareBuffer_sbuf_p1_rdat_335 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_336 = {_zz_shareBuffer_sbuf_p1_rdat_337,_zz_shareBuffer_sbuf_p1_rdat_338};
  assign _zz_shareBuffer_sbuf_p1_rdat_448 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_449 = {_zz_shareBuffer_sbuf_p1_rdat_450,_zz_shareBuffer_sbuf_p1_rdat_451};
  assign _zz_shareBuffer_sbuf_p1_rdat_561 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_562 = {_zz_shareBuffer_sbuf_p1_rdat_563,_zz_shareBuffer_sbuf_p1_rdat_564};
  assign _zz_shareBuffer_sbuf_p1_rdat_674 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_675 = {_zz_shareBuffer_sbuf_p1_rdat_676,_zz_shareBuffer_sbuf_p1_rdat_677};
  assign _zz_shareBuffer_sbuf_p1_rdat_787 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_788 = {_zz_shareBuffer_sbuf_p1_rdat_789,_zz_shareBuffer_sbuf_p1_rdat_790};
  assign _zz_shareBuffer_sbuf_p1_rdat_902 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_903 = {_zz_shareBuffer_sbuf_p1_rdat_904,_zz_shareBuffer_sbuf_p1_rdat_905};
  assign _zz_shareBuffer_sbuf_p1_rdat_1015 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1016 = {_zz_shareBuffer_sbuf_p1_rdat_1017,_zz_shareBuffer_sbuf_p1_rdat_1018};
  assign _zz_shareBuffer_sbuf_p1_rdat_1129 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1130 = {_zz_shareBuffer_sbuf_p1_rdat_1131,_zz_shareBuffer_sbuf_p1_rdat_1132};
  assign _zz_shareBuffer_sbuf_p1_rdat_1242 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1243 = {_zz_shareBuffer_sbuf_p1_rdat_1244,_zz_shareBuffer_sbuf_p1_rdat_1245};
  assign _zz_shareBuffer_sbuf_p1_rdat_1355 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1356 = {_zz_shareBuffer_sbuf_p1_rdat_1357,_zz_shareBuffer_sbuf_p1_rdat_1358};
  assign _zz_shareBuffer_sbuf_p1_rdat_1467 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1468 = {_zz_shareBuffer_sbuf_p1_rdat_1469,_zz_shareBuffer_sbuf_p1_rdat_1470};
  assign _zz_shareBuffer_sbuf_p1_rdat_1579 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1580 = {_zz_shareBuffer_sbuf_p1_rdat_1581,_zz_shareBuffer_sbuf_p1_rdat_1582};
  assign _zz_shareBuffer_sbuf_p1_rdat_1689 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1690 = {_zz_shareBuffer_sbuf_p1_rdat_1691,_zz_shareBuffer_sbuf_p1_rdat_1692};
  assign _zz_shareBuffer_sbuf_p1_rdat_6 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_7 = {_zz_shareBuffer_sbuf_p1_rdat_8,_zz_shareBuffer_sbuf_p1_rdat_9};
  assign _zz_shareBuffer_sbuf_p1_rdat_115 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_116 = {_zz_shareBuffer_sbuf_p1_rdat_117,_zz_shareBuffer_sbuf_p1_rdat_118};
  assign _zz_shareBuffer_sbuf_p1_rdat_226 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_227 = {_zz_shareBuffer_sbuf_p1_rdat_228,_zz_shareBuffer_sbuf_p1_rdat_229};
  assign _zz_shareBuffer_sbuf_p1_rdat_337 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_338 = {_zz_shareBuffer_sbuf_p1_rdat_339,_zz_shareBuffer_sbuf_p1_rdat_340};
  assign _zz_shareBuffer_sbuf_p1_rdat_450 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_451 = {_zz_shareBuffer_sbuf_p1_rdat_452,_zz_shareBuffer_sbuf_p1_rdat_453};
  assign _zz_shareBuffer_sbuf_p1_rdat_563 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_564 = {_zz_shareBuffer_sbuf_p1_rdat_565,_zz_shareBuffer_sbuf_p1_rdat_566};
  assign _zz_shareBuffer_sbuf_p1_rdat_676 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_677 = {_zz_shareBuffer_sbuf_p1_rdat_678,_zz_shareBuffer_sbuf_p1_rdat_679};
  assign _zz_shareBuffer_sbuf_p1_rdat_789 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_790 = {_zz_shareBuffer_sbuf_p1_rdat_791,_zz_shareBuffer_sbuf_p1_rdat_792};
  assign _zz_shareBuffer_sbuf_p1_rdat_904 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_905 = {_zz_shareBuffer_sbuf_p1_rdat_906,_zz_shareBuffer_sbuf_p1_rdat_907};
  assign _zz_shareBuffer_sbuf_p1_rdat_1017 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1018 = {_zz_shareBuffer_sbuf_p1_rdat_1019,_zz_shareBuffer_sbuf_p1_rdat_1020};
  assign _zz_shareBuffer_sbuf_p1_rdat_1131 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1132 = {_zz_shareBuffer_sbuf_p1_rdat_1133,_zz_shareBuffer_sbuf_p1_rdat_1134};
  assign _zz_shareBuffer_sbuf_p1_rdat_1244 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1245 = {_zz_shareBuffer_sbuf_p1_rdat_1246,_zz_shareBuffer_sbuf_p1_rdat_1247};
  assign _zz_shareBuffer_sbuf_p1_rdat_1357 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1358 = {_zz_shareBuffer_sbuf_p1_rdat_1359,_zz_shareBuffer_sbuf_p1_rdat_1360};
  assign _zz_shareBuffer_sbuf_p1_rdat_1469 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1470 = {_zz_shareBuffer_sbuf_p1_rdat_1471,_zz_shareBuffer_sbuf_p1_rdat_1472};
  assign _zz_shareBuffer_sbuf_p1_rdat_1581 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1582 = {_zz_shareBuffer_sbuf_p1_rdat_1583,_zz_shareBuffer_sbuf_p1_rdat_1584};
  assign _zz_shareBuffer_sbuf_p1_rdat_1691 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1692 = {_zz_shareBuffer_sbuf_p1_rdat_1693,_zz_shareBuffer_sbuf_p1_rdat_1694};
  assign _zz_shareBuffer_sbuf_p1_rdat_8 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_9 = {_zz_shareBuffer_sbuf_p1_rdat_10,_zz_shareBuffer_sbuf_p1_rdat_11};
  assign _zz_shareBuffer_sbuf_p1_rdat_117 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_118 = {_zz_shareBuffer_sbuf_p1_rdat_119,_zz_shareBuffer_sbuf_p1_rdat_120};
  assign _zz_shareBuffer_sbuf_p1_rdat_228 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_229 = {_zz_shareBuffer_sbuf_p1_rdat_230,_zz_shareBuffer_sbuf_p1_rdat_231};
  assign _zz_shareBuffer_sbuf_p1_rdat_339 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_340 = {_zz_shareBuffer_sbuf_p1_rdat_341,_zz_shareBuffer_sbuf_p1_rdat_342};
  assign _zz_shareBuffer_sbuf_p1_rdat_452 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_453 = {_zz_shareBuffer_sbuf_p1_rdat_454,_zz_shareBuffer_sbuf_p1_rdat_455};
  assign _zz_shareBuffer_sbuf_p1_rdat_565 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_566 = {_zz_shareBuffer_sbuf_p1_rdat_567,_zz_shareBuffer_sbuf_p1_rdat_568};
  assign _zz_shareBuffer_sbuf_p1_rdat_678 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_679 = {_zz_shareBuffer_sbuf_p1_rdat_680,_zz_shareBuffer_sbuf_p1_rdat_681};
  assign _zz_shareBuffer_sbuf_p1_rdat_791 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_792 = {_zz_shareBuffer_sbuf_p1_rdat_793,_zz_shareBuffer_sbuf_p1_rdat_794};
  assign _zz_shareBuffer_sbuf_p1_rdat_906 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_907 = {_zz_shareBuffer_sbuf_p1_rdat_908,_zz_shareBuffer_sbuf_p1_rdat_909};
  assign _zz_shareBuffer_sbuf_p1_rdat_1019 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1020 = {_zz_shareBuffer_sbuf_p1_rdat_1021,_zz_shareBuffer_sbuf_p1_rdat_1022};
  assign _zz_shareBuffer_sbuf_p1_rdat_1133 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1134 = {_zz_shareBuffer_sbuf_p1_rdat_1135,_zz_shareBuffer_sbuf_p1_rdat_1136};
  assign _zz_shareBuffer_sbuf_p1_rdat_1246 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1247 = {_zz_shareBuffer_sbuf_p1_rdat_1248,_zz_shareBuffer_sbuf_p1_rdat_1249};
  assign _zz_shareBuffer_sbuf_p1_rdat_1359 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1360 = {_zz_shareBuffer_sbuf_p1_rdat_1361,_zz_shareBuffer_sbuf_p1_rdat_1362};
  assign _zz_shareBuffer_sbuf_p1_rdat_1471 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1472 = {_zz_shareBuffer_sbuf_p1_rdat_1473,_zz_shareBuffer_sbuf_p1_rdat_1474};
  assign _zz_shareBuffer_sbuf_p1_rdat_1583 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1584 = {_zz_shareBuffer_sbuf_p1_rdat_1585,_zz_shareBuffer_sbuf_p1_rdat_1586};
  assign _zz_shareBuffer_sbuf_p1_rdat_1693 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1694 = {_zz_shareBuffer_sbuf_p1_rdat_1695,_zz_shareBuffer_sbuf_p1_rdat_1696};
  assign _zz_shareBuffer_sbuf_p1_rdat_10 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_11 = {_zz_shareBuffer_sbuf_p1_rdat_12,_zz_shareBuffer_sbuf_p1_rdat_13};
  assign _zz_shareBuffer_sbuf_p1_rdat_119 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_120 = {_zz_shareBuffer_sbuf_p1_rdat_121,_zz_shareBuffer_sbuf_p1_rdat_122};
  assign _zz_shareBuffer_sbuf_p1_rdat_230 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_231 = {_zz_shareBuffer_sbuf_p1_rdat_232,_zz_shareBuffer_sbuf_p1_rdat_233};
  assign _zz_shareBuffer_sbuf_p1_rdat_341 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_342 = {_zz_shareBuffer_sbuf_p1_rdat_343,_zz_shareBuffer_sbuf_p1_rdat_344};
  assign _zz_shareBuffer_sbuf_p1_rdat_454 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_455 = {_zz_shareBuffer_sbuf_p1_rdat_456,_zz_shareBuffer_sbuf_p1_rdat_457};
  assign _zz_shareBuffer_sbuf_p1_rdat_567 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_568 = {_zz_shareBuffer_sbuf_p1_rdat_569,_zz_shareBuffer_sbuf_p1_rdat_570};
  assign _zz_shareBuffer_sbuf_p1_rdat_680 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_681 = {_zz_shareBuffer_sbuf_p1_rdat_682,_zz_shareBuffer_sbuf_p1_rdat_683};
  assign _zz_shareBuffer_sbuf_p1_rdat_793 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_794 = {_zz_shareBuffer_sbuf_p1_rdat_795,_zz_shareBuffer_sbuf_p1_rdat_796};
  assign _zz_shareBuffer_sbuf_p1_rdat_908 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_909 = {_zz_shareBuffer_sbuf_p1_rdat_910,_zz_shareBuffer_sbuf_p1_rdat_911};
  assign _zz_shareBuffer_sbuf_p1_rdat_1021 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1022 = {_zz_shareBuffer_sbuf_p1_rdat_1023,_zz_shareBuffer_sbuf_p1_rdat_1024};
  assign _zz_shareBuffer_sbuf_p1_rdat_1135 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1136 = {_zz_shareBuffer_sbuf_p1_rdat_1137,_zz_shareBuffer_sbuf_p1_rdat_1138};
  assign _zz_shareBuffer_sbuf_p1_rdat_1248 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1249 = {_zz_shareBuffer_sbuf_p1_rdat_1250,_zz_shareBuffer_sbuf_p1_rdat_1251};
  assign _zz_shareBuffer_sbuf_p1_rdat_1361 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1362 = {_zz_shareBuffer_sbuf_p1_rdat_1363,_zz_shareBuffer_sbuf_p1_rdat_1364};
  assign _zz_shareBuffer_sbuf_p1_rdat_1473 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1474 = {_zz_shareBuffer_sbuf_p1_rdat_1475,_zz_shareBuffer_sbuf_p1_rdat_1476};
  assign _zz_shareBuffer_sbuf_p1_rdat_1585 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1586 = {_zz_shareBuffer_sbuf_p1_rdat_1587,_zz_shareBuffer_sbuf_p1_rdat_1588};
  assign _zz_shareBuffer_sbuf_p1_rdat_1695 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1696 = {_zz_shareBuffer_sbuf_p1_rdat_1697,_zz_shareBuffer_sbuf_p1_rdat_1698};
  assign _zz_shareBuffer_sbuf_p1_rdat_12 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_13 = {_zz_shareBuffer_sbuf_p1_rdat_14,_zz_shareBuffer_sbuf_p1_rdat_15};
  assign _zz_shareBuffer_sbuf_p1_rdat_121 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_122 = {_zz_shareBuffer_sbuf_p1_rdat_123,_zz_shareBuffer_sbuf_p1_rdat_124};
  assign _zz_shareBuffer_sbuf_p1_rdat_232 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_233 = {_zz_shareBuffer_sbuf_p1_rdat_234,_zz_shareBuffer_sbuf_p1_rdat_235};
  assign _zz_shareBuffer_sbuf_p1_rdat_343 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_344 = {_zz_shareBuffer_sbuf_p1_rdat_345,_zz_shareBuffer_sbuf_p1_rdat_346};
  assign _zz_shareBuffer_sbuf_p1_rdat_456 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_457 = {_zz_shareBuffer_sbuf_p1_rdat_458,_zz_shareBuffer_sbuf_p1_rdat_459};
  assign _zz_shareBuffer_sbuf_p1_rdat_569 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_570 = {_zz_shareBuffer_sbuf_p1_rdat_571,_zz_shareBuffer_sbuf_p1_rdat_572};
  assign _zz_shareBuffer_sbuf_p1_rdat_682 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_683 = {_zz_shareBuffer_sbuf_p1_rdat_684,_zz_shareBuffer_sbuf_p1_rdat_685};
  assign _zz_shareBuffer_sbuf_p1_rdat_795 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_796 = {_zz_shareBuffer_sbuf_p1_rdat_797,_zz_shareBuffer_sbuf_p1_rdat_798};
  assign _zz_shareBuffer_sbuf_p1_rdat_910 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_911 = {_zz_shareBuffer_sbuf_p1_rdat_912,_zz_shareBuffer_sbuf_p1_rdat_913};
  assign _zz_shareBuffer_sbuf_p1_rdat_1023 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1024 = {_zz_shareBuffer_sbuf_p1_rdat_1025,_zz_shareBuffer_sbuf_p1_rdat_1026};
  assign _zz_shareBuffer_sbuf_p1_rdat_1137 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1138 = {_zz_shareBuffer_sbuf_p1_rdat_1139,_zz_shareBuffer_sbuf_p1_rdat_1140};
  assign _zz_shareBuffer_sbuf_p1_rdat_1250 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1251 = {_zz_shareBuffer_sbuf_p1_rdat_1252,_zz_shareBuffer_sbuf_p1_rdat_1253};
  assign _zz_shareBuffer_sbuf_p1_rdat_1363 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1364 = {_zz_shareBuffer_sbuf_p1_rdat_1365,_zz_shareBuffer_sbuf_p1_rdat_1366};
  assign _zz_shareBuffer_sbuf_p1_rdat_1475 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1476 = {_zz_shareBuffer_sbuf_p1_rdat_1477,_zz_shareBuffer_sbuf_p1_rdat_1478};
  assign _zz_shareBuffer_sbuf_p1_rdat_1587 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1588 = {_zz_shareBuffer_sbuf_p1_rdat_1589,_zz_shareBuffer_sbuf_p1_rdat_1590};
  assign _zz_shareBuffer_sbuf_p1_rdat_1697 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1698 = {_zz_shareBuffer_sbuf_p1_rdat_1699,_zz_shareBuffer_sbuf_p1_rdat_1700};
  assign _zz_shareBuffer_sbuf_p1_rdat_14 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_15 = {_zz_shareBuffer_sbuf_p1_rdat_16,_zz_shareBuffer_sbuf_p1_rdat_17};
  assign _zz_shareBuffer_sbuf_p1_rdat_123 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_124 = {_zz_shareBuffer_sbuf_p1_rdat_125,_zz_shareBuffer_sbuf_p1_rdat_126};
  assign _zz_shareBuffer_sbuf_p1_rdat_234 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_235 = {_zz_shareBuffer_sbuf_p1_rdat_236,_zz_shareBuffer_sbuf_p1_rdat_237};
  assign _zz_shareBuffer_sbuf_p1_rdat_345 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_346 = {_zz_shareBuffer_sbuf_p1_rdat_347,_zz_shareBuffer_sbuf_p1_rdat_348};
  assign _zz_shareBuffer_sbuf_p1_rdat_458 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_459 = {_zz_shareBuffer_sbuf_p1_rdat_460,_zz_shareBuffer_sbuf_p1_rdat_461};
  assign _zz_shareBuffer_sbuf_p1_rdat_571 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_572 = {_zz_shareBuffer_sbuf_p1_rdat_573,_zz_shareBuffer_sbuf_p1_rdat_574};
  assign _zz_shareBuffer_sbuf_p1_rdat_684 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_685 = {_zz_shareBuffer_sbuf_p1_rdat_686,_zz_shareBuffer_sbuf_p1_rdat_687};
  assign _zz_shareBuffer_sbuf_p1_rdat_797 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_798 = {_zz_shareBuffer_sbuf_p1_rdat_799,_zz_shareBuffer_sbuf_p1_rdat_800};
  assign _zz_shareBuffer_sbuf_p1_rdat_912 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_913 = {_zz_shareBuffer_sbuf_p1_rdat_914,_zz_shareBuffer_sbuf_p1_rdat_915};
  assign _zz_shareBuffer_sbuf_p1_rdat_1025 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1026 = {_zz_shareBuffer_sbuf_p1_rdat_1027,_zz_shareBuffer_sbuf_p1_rdat_1028};
  assign _zz_shareBuffer_sbuf_p1_rdat_1139 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1140 = {_zz_shareBuffer_sbuf_p1_rdat_1141,_zz_shareBuffer_sbuf_p1_rdat_1142};
  assign _zz_shareBuffer_sbuf_p1_rdat_1252 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1253 = {_zz_shareBuffer_sbuf_p1_rdat_1254,_zz_shareBuffer_sbuf_p1_rdat_1255};
  assign _zz_shareBuffer_sbuf_p1_rdat_1365 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1366 = {_zz_shareBuffer_sbuf_p1_rdat_1367,_zz_shareBuffer_sbuf_p1_rdat_1368};
  assign _zz_shareBuffer_sbuf_p1_rdat_1477 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1478 = {_zz_shareBuffer_sbuf_p1_rdat_1479,_zz_shareBuffer_sbuf_p1_rdat_1480};
  assign _zz_shareBuffer_sbuf_p1_rdat_1589 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1590 = {_zz_shareBuffer_sbuf_p1_rdat_1591,_zz_shareBuffer_sbuf_p1_rdat_1592};
  assign _zz_shareBuffer_sbuf_p1_rdat_1699 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1700 = {_zz_shareBuffer_sbuf_p1_rdat_1701,_zz_shareBuffer_sbuf_p1_rdat_1702};
  assign _zz_shareBuffer_sbuf_p1_rdat_16 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_17 = {_zz_shareBuffer_sbuf_p1_rdat_18,_zz_shareBuffer_sbuf_p1_rdat_19};
  assign _zz_shareBuffer_sbuf_p1_rdat_125 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_126 = {_zz_shareBuffer_sbuf_p1_rdat_127,_zz_shareBuffer_sbuf_p1_rdat_128};
  assign _zz_shareBuffer_sbuf_p1_rdat_236 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_237 = {_zz_shareBuffer_sbuf_p1_rdat_238,_zz_shareBuffer_sbuf_p1_rdat_239};
  assign _zz_shareBuffer_sbuf_p1_rdat_347 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_348 = {_zz_shareBuffer_sbuf_p1_rdat_349,_zz_shareBuffer_sbuf_p1_rdat_350};
  assign _zz_shareBuffer_sbuf_p1_rdat_460 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_461 = {_zz_shareBuffer_sbuf_p1_rdat_462,_zz_shareBuffer_sbuf_p1_rdat_463};
  assign _zz_shareBuffer_sbuf_p1_rdat_573 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_574 = {_zz_shareBuffer_sbuf_p1_rdat_575,_zz_shareBuffer_sbuf_p1_rdat_576};
  assign _zz_shareBuffer_sbuf_p1_rdat_686 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_687 = {_zz_shareBuffer_sbuf_p1_rdat_688,_zz_shareBuffer_sbuf_p1_rdat_689};
  assign _zz_shareBuffer_sbuf_p1_rdat_799 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_800 = {_zz_shareBuffer_sbuf_p1_rdat_801,_zz_shareBuffer_sbuf_p1_rdat_802};
  assign _zz_shareBuffer_sbuf_p1_rdat_914 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_915 = {_zz_shareBuffer_sbuf_p1_rdat_916,_zz_shareBuffer_sbuf_p1_rdat_917};
  assign _zz_shareBuffer_sbuf_p1_rdat_1027 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1028 = {_zz_shareBuffer_sbuf_p1_rdat_1029,_zz_shareBuffer_sbuf_p1_rdat_1030};
  assign _zz_shareBuffer_sbuf_p1_rdat_1141 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1142 = {_zz_shareBuffer_sbuf_p1_rdat_1143,_zz_shareBuffer_sbuf_p1_rdat_1144};
  assign _zz_shareBuffer_sbuf_p1_rdat_1254 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1255 = {_zz_shareBuffer_sbuf_p1_rdat_1256,_zz_shareBuffer_sbuf_p1_rdat_1257};
  assign _zz_shareBuffer_sbuf_p1_rdat_1367 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1368 = {_zz_shareBuffer_sbuf_p1_rdat_1369,_zz_shareBuffer_sbuf_p1_rdat_1370};
  assign _zz_shareBuffer_sbuf_p1_rdat_1479 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1480 = {_zz_shareBuffer_sbuf_p1_rdat_1481,_zz_shareBuffer_sbuf_p1_rdat_1482};
  assign _zz_shareBuffer_sbuf_p1_rdat_1591 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1592 = {_zz_shareBuffer_sbuf_p1_rdat_1593,_zz_shareBuffer_sbuf_p1_rdat_1594};
  assign _zz_shareBuffer_sbuf_p1_rdat_1701 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1702 = {_zz_shareBuffer_sbuf_p1_rdat_1703,_zz_shareBuffer_sbuf_p1_rdat_1704};
  assign _zz_shareBuffer_sbuf_p1_rdat_18 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_19 = {_zz_shareBuffer_sbuf_p1_rdat_20,_zz_shareBuffer_sbuf_p1_rdat_21};
  assign _zz_shareBuffer_sbuf_p1_rdat_127 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_128 = {_zz_shareBuffer_sbuf_p1_rdat_129,_zz_shareBuffer_sbuf_p1_rdat_130};
  assign _zz_shareBuffer_sbuf_p1_rdat_238 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_239 = {_zz_shareBuffer_sbuf_p1_rdat_240,_zz_shareBuffer_sbuf_p1_rdat_241};
  assign _zz_shareBuffer_sbuf_p1_rdat_349 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_350 = {_zz_shareBuffer_sbuf_p1_rdat_351,_zz_shareBuffer_sbuf_p1_rdat_352};
  assign _zz_shareBuffer_sbuf_p1_rdat_462 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_463 = {_zz_shareBuffer_sbuf_p1_rdat_464,_zz_shareBuffer_sbuf_p1_rdat_465};
  assign _zz_shareBuffer_sbuf_p1_rdat_575 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_576 = {_zz_shareBuffer_sbuf_p1_rdat_577,_zz_shareBuffer_sbuf_p1_rdat_578};
  assign _zz_shareBuffer_sbuf_p1_rdat_688 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_689 = {_zz_shareBuffer_sbuf_p1_rdat_690,_zz_shareBuffer_sbuf_p1_rdat_691};
  assign _zz_shareBuffer_sbuf_p1_rdat_801 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_802 = {_zz_shareBuffer_sbuf_p1_rdat_803,_zz_shareBuffer_sbuf_p1_rdat_804};
  assign _zz_shareBuffer_sbuf_p1_rdat_916 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_917 = {_zz_shareBuffer_sbuf_p1_rdat_918,_zz_shareBuffer_sbuf_p1_rdat_919};
  assign _zz_shareBuffer_sbuf_p1_rdat_1029 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1030 = {_zz_shareBuffer_sbuf_p1_rdat_1031,_zz_shareBuffer_sbuf_p1_rdat_1032};
  assign _zz_shareBuffer_sbuf_p1_rdat_1143 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1144 = {_zz_shareBuffer_sbuf_p1_rdat_1145,_zz_shareBuffer_sbuf_p1_rdat_1146};
  assign _zz_shareBuffer_sbuf_p1_rdat_1256 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1257 = {_zz_shareBuffer_sbuf_p1_rdat_1258,_zz_shareBuffer_sbuf_p1_rdat_1259};
  assign _zz_shareBuffer_sbuf_p1_rdat_1369 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1370 = {_zz_shareBuffer_sbuf_p1_rdat_1371,_zz_shareBuffer_sbuf_p1_rdat_1372};
  assign _zz_shareBuffer_sbuf_p1_rdat_1481 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1482 = {_zz_shareBuffer_sbuf_p1_rdat_1483,_zz_shareBuffer_sbuf_p1_rdat_1484};
  assign _zz_shareBuffer_sbuf_p1_rdat_1593 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1594 = {_zz_shareBuffer_sbuf_p1_rdat_1595,_zz_shareBuffer_sbuf_p1_rdat_1596};
  assign _zz_shareBuffer_sbuf_p1_rdat_1703 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1704 = {_zz_shareBuffer_sbuf_p1_rdat_1705,_zz_shareBuffer_sbuf_p1_rdat_1706};
  assign _zz_shareBuffer_sbuf_p1_rdat_20 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_21 = {_zz_shareBuffer_sbuf_p1_rdat_22,_zz_shareBuffer_sbuf_p1_rdat_23};
  assign _zz_shareBuffer_sbuf_p1_rdat_129 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_130 = {_zz_shareBuffer_sbuf_p1_rdat_131,_zz_shareBuffer_sbuf_p1_rdat_132};
  assign _zz_shareBuffer_sbuf_p1_rdat_240 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_241 = {_zz_shareBuffer_sbuf_p1_rdat_242,_zz_shareBuffer_sbuf_p1_rdat_243};
  assign _zz_shareBuffer_sbuf_p1_rdat_351 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_352 = {_zz_shareBuffer_sbuf_p1_rdat_353,_zz_shareBuffer_sbuf_p1_rdat_354};
  assign _zz_shareBuffer_sbuf_p1_rdat_464 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_465 = {_zz_shareBuffer_sbuf_p1_rdat_466,_zz_shareBuffer_sbuf_p1_rdat_467};
  assign _zz_shareBuffer_sbuf_p1_rdat_577 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_578 = {_zz_shareBuffer_sbuf_p1_rdat_579,_zz_shareBuffer_sbuf_p1_rdat_580};
  assign _zz_shareBuffer_sbuf_p1_rdat_690 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_691 = {_zz_shareBuffer_sbuf_p1_rdat_692,_zz_shareBuffer_sbuf_p1_rdat_693};
  assign _zz_shareBuffer_sbuf_p1_rdat_803 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_804 = {_zz_shareBuffer_sbuf_p1_rdat_805,_zz_shareBuffer_sbuf_p1_rdat_806};
  assign _zz_shareBuffer_sbuf_p1_rdat_918 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_919 = {_zz_shareBuffer_sbuf_p1_rdat_920,_zz_shareBuffer_sbuf_p1_rdat_921};
  assign _zz_shareBuffer_sbuf_p1_rdat_1031 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1032 = {_zz_shareBuffer_sbuf_p1_rdat_1033,_zz_shareBuffer_sbuf_p1_rdat_1034};
  assign _zz_shareBuffer_sbuf_p1_rdat_1145 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1146 = {_zz_shareBuffer_sbuf_p1_rdat_1147,_zz_shareBuffer_sbuf_p1_rdat_1148};
  assign _zz_shareBuffer_sbuf_p1_rdat_1258 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1259 = {_zz_shareBuffer_sbuf_p1_rdat_1260,_zz_shareBuffer_sbuf_p1_rdat_1261};
  assign _zz_shareBuffer_sbuf_p1_rdat_1371 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1372 = {_zz_shareBuffer_sbuf_p1_rdat_1373,_zz_shareBuffer_sbuf_p1_rdat_1374};
  assign _zz_shareBuffer_sbuf_p1_rdat_1483 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1484 = {_zz_shareBuffer_sbuf_p1_rdat_1485,_zz_shareBuffer_sbuf_p1_rdat_1486};
  assign _zz_shareBuffer_sbuf_p1_rdat_1595 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1596 = {_zz_shareBuffer_sbuf_p1_rdat_1597,_zz_shareBuffer_sbuf_p1_rdat_1598};
  assign _zz_shareBuffer_sbuf_p1_rdat_1705 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1706 = {_zz_shareBuffer_sbuf_p1_rdat_1707,_zz_shareBuffer_sbuf_p1_rdat_1708};
  assign _zz_shareBuffer_sbuf_p1_rdat_22 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_23 = {_zz_shareBuffer_sbuf_p1_rdat_24,_zz_shareBuffer_sbuf_p1_rdat_25};
  assign _zz_shareBuffer_sbuf_p1_rdat_131 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_132 = {_zz_shareBuffer_sbuf_p1_rdat_133,_zz_shareBuffer_sbuf_p1_rdat_134};
  assign _zz_shareBuffer_sbuf_p1_rdat_242 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_243 = {_zz_shareBuffer_sbuf_p1_rdat_244,_zz_shareBuffer_sbuf_p1_rdat_245};
  assign _zz_shareBuffer_sbuf_p1_rdat_353 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_354 = {_zz_shareBuffer_sbuf_p1_rdat_355,_zz_shareBuffer_sbuf_p1_rdat_356};
  assign _zz_shareBuffer_sbuf_p1_rdat_466 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_467 = {_zz_shareBuffer_sbuf_p1_rdat_468,_zz_shareBuffer_sbuf_p1_rdat_469};
  assign _zz_shareBuffer_sbuf_p1_rdat_579 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_580 = {_zz_shareBuffer_sbuf_p1_rdat_581,_zz_shareBuffer_sbuf_p1_rdat_582};
  assign _zz_shareBuffer_sbuf_p1_rdat_692 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_693 = {_zz_shareBuffer_sbuf_p1_rdat_694,_zz_shareBuffer_sbuf_p1_rdat_695};
  assign _zz_shareBuffer_sbuf_p1_rdat_805 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_806 = {_zz_shareBuffer_sbuf_p1_rdat_807,_zz_shareBuffer_sbuf_p1_rdat_808};
  assign _zz_shareBuffer_sbuf_p1_rdat_920 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_921 = {_zz_shareBuffer_sbuf_p1_rdat_922,_zz_shareBuffer_sbuf_p1_rdat_923};
  assign _zz_shareBuffer_sbuf_p1_rdat_1033 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1034 = {_zz_shareBuffer_sbuf_p1_rdat_1035,_zz_shareBuffer_sbuf_p1_rdat_1036};
  assign _zz_shareBuffer_sbuf_p1_rdat_1147 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1148 = {_zz_shareBuffer_sbuf_p1_rdat_1149,_zz_shareBuffer_sbuf_p1_rdat_1150};
  assign _zz_shareBuffer_sbuf_p1_rdat_1260 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1261 = {_zz_shareBuffer_sbuf_p1_rdat_1262,_zz_shareBuffer_sbuf_p1_rdat_1263};
  assign _zz_shareBuffer_sbuf_p1_rdat_1373 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1374 = {_zz_shareBuffer_sbuf_p1_rdat_1375,_zz_shareBuffer_sbuf_p1_rdat_1376};
  assign _zz_shareBuffer_sbuf_p1_rdat_1485 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1486 = {_zz_shareBuffer_sbuf_p1_rdat_1487,_zz_shareBuffer_sbuf_p1_rdat_1488};
  assign _zz_shareBuffer_sbuf_p1_rdat_1597 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1598 = {_zz_shareBuffer_sbuf_p1_rdat_1599,_zz_shareBuffer_sbuf_p1_rdat_1600};
  assign _zz_shareBuffer_sbuf_p1_rdat_1707 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1708 = {_zz_shareBuffer_sbuf_p1_rdat_1709,_zz_shareBuffer_sbuf_p1_rdat_1710};
  assign _zz_shareBuffer_sbuf_p1_rdat_24 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_25 = {_zz_shareBuffer_sbuf_p1_rdat_26,_zz_shareBuffer_sbuf_p1_rdat_27};
  assign _zz_shareBuffer_sbuf_p1_rdat_133 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_134 = {_zz_shareBuffer_sbuf_p1_rdat_135,_zz_shareBuffer_sbuf_p1_rdat_136};
  assign _zz_shareBuffer_sbuf_p1_rdat_244 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_245 = {_zz_shareBuffer_sbuf_p1_rdat_246,_zz_shareBuffer_sbuf_p1_rdat_247};
  assign _zz_shareBuffer_sbuf_p1_rdat_355 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_356 = {_zz_shareBuffer_sbuf_p1_rdat_357,_zz_shareBuffer_sbuf_p1_rdat_358};
  assign _zz_shareBuffer_sbuf_p1_rdat_468 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_469 = {_zz_shareBuffer_sbuf_p1_rdat_470,_zz_shareBuffer_sbuf_p1_rdat_471};
  assign _zz_shareBuffer_sbuf_p1_rdat_581 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_582 = {_zz_shareBuffer_sbuf_p1_rdat_583,_zz_shareBuffer_sbuf_p1_rdat_584};
  assign _zz_shareBuffer_sbuf_p1_rdat_694 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_695 = {_zz_shareBuffer_sbuf_p1_rdat_696,_zz_shareBuffer_sbuf_p1_rdat_697};
  assign _zz_shareBuffer_sbuf_p1_rdat_807 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_808 = {_zz_shareBuffer_sbuf_p1_rdat_809,_zz_shareBuffer_sbuf_p1_rdat_810};
  assign _zz_shareBuffer_sbuf_p1_rdat_922 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_923 = {_zz_shareBuffer_sbuf_p1_rdat_924,_zz_shareBuffer_sbuf_p1_rdat_925};
  assign _zz_shareBuffer_sbuf_p1_rdat_1035 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1036 = {_zz_shareBuffer_sbuf_p1_rdat_1037,_zz_shareBuffer_sbuf_p1_rdat_1038};
  assign _zz_shareBuffer_sbuf_p1_rdat_1149 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1150 = {_zz_shareBuffer_sbuf_p1_rdat_1151,_zz_shareBuffer_sbuf_p1_rdat_1152};
  assign _zz_shareBuffer_sbuf_p1_rdat_1262 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1263 = {_zz_shareBuffer_sbuf_p1_rdat_1264,_zz_shareBuffer_sbuf_p1_rdat_1265};
  assign _zz_shareBuffer_sbuf_p1_rdat_1375 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1376 = {_zz_shareBuffer_sbuf_p1_rdat_1377,_zz_shareBuffer_sbuf_p1_rdat_1378};
  assign _zz_shareBuffer_sbuf_p1_rdat_1487 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1488 = {_zz_shareBuffer_sbuf_p1_rdat_1489,_zz_shareBuffer_sbuf_p1_rdat_1490};
  assign _zz_shareBuffer_sbuf_p1_rdat_1599 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1600 = {_zz_shareBuffer_sbuf_p1_rdat_1601,_zz_shareBuffer_sbuf_p1_rdat_1602};
  assign _zz_shareBuffer_sbuf_p1_rdat_1709 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1710 = {_zz_shareBuffer_sbuf_p1_rdat_1711,_zz_shareBuffer_sbuf_p1_rdat_1712};
  assign _zz_shareBuffer_sbuf_p1_rdat_26 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_27 = {_zz_shareBuffer_sbuf_p1_rdat_28,_zz_shareBuffer_sbuf_p1_rdat_29};
  assign _zz_shareBuffer_sbuf_p1_rdat_135 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_136 = {_zz_shareBuffer_sbuf_p1_rdat_137,_zz_shareBuffer_sbuf_p1_rdat_138};
  assign _zz_shareBuffer_sbuf_p1_rdat_246 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_247 = {_zz_shareBuffer_sbuf_p1_rdat_248,_zz_shareBuffer_sbuf_p1_rdat_249};
  assign _zz_shareBuffer_sbuf_p1_rdat_357 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_358 = {_zz_shareBuffer_sbuf_p1_rdat_359,_zz_shareBuffer_sbuf_p1_rdat_360};
  assign _zz_shareBuffer_sbuf_p1_rdat_470 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_471 = {_zz_shareBuffer_sbuf_p1_rdat_472,_zz_shareBuffer_sbuf_p1_rdat_473};
  assign _zz_shareBuffer_sbuf_p1_rdat_583 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_584 = {_zz_shareBuffer_sbuf_p1_rdat_585,_zz_shareBuffer_sbuf_p1_rdat_586};
  assign _zz_shareBuffer_sbuf_p1_rdat_696 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_697 = {_zz_shareBuffer_sbuf_p1_rdat_698,_zz_shareBuffer_sbuf_p1_rdat_699};
  assign _zz_shareBuffer_sbuf_p1_rdat_809 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_810 = {_zz_shareBuffer_sbuf_p1_rdat_811,_zz_shareBuffer_sbuf_p1_rdat_812};
  assign _zz_shareBuffer_sbuf_p1_rdat_924 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_925 = {_zz_shareBuffer_sbuf_p1_rdat_926,_zz_shareBuffer_sbuf_p1_rdat_927};
  assign _zz_shareBuffer_sbuf_p1_rdat_1037 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1038 = {_zz_shareBuffer_sbuf_p1_rdat_1039,_zz_shareBuffer_sbuf_p1_rdat_1040};
  assign _zz_shareBuffer_sbuf_p1_rdat_1151 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1152 = {_zz_shareBuffer_sbuf_p1_rdat_1153,_zz_shareBuffer_sbuf_p1_rdat_1154};
  assign _zz_shareBuffer_sbuf_p1_rdat_1264 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1265 = {_zz_shareBuffer_sbuf_p1_rdat_1266,_zz_shareBuffer_sbuf_p1_rdat_1267};
  assign _zz_shareBuffer_sbuf_p1_rdat_1377 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1378 = {_zz_shareBuffer_sbuf_p1_rdat_1379,_zz_shareBuffer_sbuf_p1_rdat_1380};
  assign _zz_shareBuffer_sbuf_p1_rdat_1489 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1490 = {_zz_shareBuffer_sbuf_p1_rdat_1491,_zz_shareBuffer_sbuf_p1_rdat_1492};
  assign _zz_shareBuffer_sbuf_p1_rdat_1601 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1602 = {_zz_shareBuffer_sbuf_p1_rdat_1603,_zz_shareBuffer_sbuf_p1_rdat_1604};
  assign _zz_shareBuffer_sbuf_p1_rdat_1711 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1712 = {_zz_shareBuffer_sbuf_p1_rdat_1713,_zz_shareBuffer_sbuf_p1_rdat_1714};
  assign _zz_shareBuffer_sbuf_p1_rdat_28 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_29 = {_zz_shareBuffer_sbuf_p1_rdat_30,_zz_shareBuffer_sbuf_p1_rdat_31};
  assign _zz_shareBuffer_sbuf_p1_rdat_137 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_138 = {_zz_shareBuffer_sbuf_p1_rdat_139,_zz_shareBuffer_sbuf_p1_rdat_140};
  assign _zz_shareBuffer_sbuf_p1_rdat_248 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_249 = {_zz_shareBuffer_sbuf_p1_rdat_250,_zz_shareBuffer_sbuf_p1_rdat_251};
  assign _zz_shareBuffer_sbuf_p1_rdat_359 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_360 = {_zz_shareBuffer_sbuf_p1_rdat_361,_zz_shareBuffer_sbuf_p1_rdat_362};
  assign _zz_shareBuffer_sbuf_p1_rdat_472 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_473 = {_zz_shareBuffer_sbuf_p1_rdat_474,_zz_shareBuffer_sbuf_p1_rdat_475};
  assign _zz_shareBuffer_sbuf_p1_rdat_585 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_586 = {_zz_shareBuffer_sbuf_p1_rdat_587,_zz_shareBuffer_sbuf_p1_rdat_588};
  assign _zz_shareBuffer_sbuf_p1_rdat_698 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_699 = {_zz_shareBuffer_sbuf_p1_rdat_700,_zz_shareBuffer_sbuf_p1_rdat_701};
  assign _zz_shareBuffer_sbuf_p1_rdat_811 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_812 = {_zz_shareBuffer_sbuf_p1_rdat_813,_zz_shareBuffer_sbuf_p1_rdat_814};
  assign _zz_shareBuffer_sbuf_p1_rdat_926 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_927 = {_zz_shareBuffer_sbuf_p1_rdat_928,_zz_shareBuffer_sbuf_p1_rdat_929};
  assign _zz_shareBuffer_sbuf_p1_rdat_1039 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1040 = {_zz_shareBuffer_sbuf_p1_rdat_1041,_zz_shareBuffer_sbuf_p1_rdat_1042};
  assign _zz_shareBuffer_sbuf_p1_rdat_1153 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1154 = {_zz_shareBuffer_sbuf_p1_rdat_1155,_zz_shareBuffer_sbuf_p1_rdat_1156};
  assign _zz_shareBuffer_sbuf_p1_rdat_1266 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1267 = {_zz_shareBuffer_sbuf_p1_rdat_1268,_zz_shareBuffer_sbuf_p1_rdat_1269};
  assign _zz_shareBuffer_sbuf_p1_rdat_1379 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1380 = {_zz_shareBuffer_sbuf_p1_rdat_1381,_zz_shareBuffer_sbuf_p1_rdat_1382};
  assign _zz_shareBuffer_sbuf_p1_rdat_1491 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1492 = {_zz_shareBuffer_sbuf_p1_rdat_1493,_zz_shareBuffer_sbuf_p1_rdat_1494};
  assign _zz_shareBuffer_sbuf_p1_rdat_1603 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1604 = {_zz_shareBuffer_sbuf_p1_rdat_1605,_zz_shareBuffer_sbuf_p1_rdat_1606};
  assign _zz_shareBuffer_sbuf_p1_rdat_1713 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1714 = {_zz_shareBuffer_sbuf_p1_rdat_1715,_zz_shareBuffer_sbuf_p1_rdat_1716};
  assign _zz_shareBuffer_sbuf_p1_rdat_30 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_31 = {_zz_shareBuffer_sbuf_p1_rdat_32,_zz_shareBuffer_sbuf_p1_rdat_33};
  assign _zz_shareBuffer_sbuf_p1_rdat_139 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_140 = {_zz_shareBuffer_sbuf_p1_rdat_141,_zz_shareBuffer_sbuf_p1_rdat_142};
  assign _zz_shareBuffer_sbuf_p1_rdat_250 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_251 = {_zz_shareBuffer_sbuf_p1_rdat_252,_zz_shareBuffer_sbuf_p1_rdat_253};
  assign _zz_shareBuffer_sbuf_p1_rdat_361 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_362 = {_zz_shareBuffer_sbuf_p1_rdat_363,_zz_shareBuffer_sbuf_p1_rdat_364};
  assign _zz_shareBuffer_sbuf_p1_rdat_474 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_475 = {_zz_shareBuffer_sbuf_p1_rdat_476,_zz_shareBuffer_sbuf_p1_rdat_477};
  assign _zz_shareBuffer_sbuf_p1_rdat_587 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_588 = {_zz_shareBuffer_sbuf_p1_rdat_589,_zz_shareBuffer_sbuf_p1_rdat_590};
  assign _zz_shareBuffer_sbuf_p1_rdat_700 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_701 = {_zz_shareBuffer_sbuf_p1_rdat_702,_zz_shareBuffer_sbuf_p1_rdat_703};
  assign _zz_shareBuffer_sbuf_p1_rdat_813 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_814 = {_zz_shareBuffer_sbuf_p1_rdat_815,_zz_shareBuffer_sbuf_p1_rdat_816};
  assign _zz_shareBuffer_sbuf_p1_rdat_928 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_929 = {_zz_shareBuffer_sbuf_p1_rdat_930,_zz_shareBuffer_sbuf_p1_rdat_931};
  assign _zz_shareBuffer_sbuf_p1_rdat_1041 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1042 = {_zz_shareBuffer_sbuf_p1_rdat_1043,_zz_shareBuffer_sbuf_p1_rdat_1044};
  assign _zz_shareBuffer_sbuf_p1_rdat_1155 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1156 = {_zz_shareBuffer_sbuf_p1_rdat_1157,_zz_shareBuffer_sbuf_p1_rdat_1158};
  assign _zz_shareBuffer_sbuf_p1_rdat_1268 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1269 = {_zz_shareBuffer_sbuf_p1_rdat_1270,_zz_shareBuffer_sbuf_p1_rdat_1271};
  assign _zz_shareBuffer_sbuf_p1_rdat_1381 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1382 = {_zz_shareBuffer_sbuf_p1_rdat_1383,_zz_shareBuffer_sbuf_p1_rdat_1384};
  assign _zz_shareBuffer_sbuf_p1_rdat_1493 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1494 = {_zz_shareBuffer_sbuf_p1_rdat_1495,_zz_shareBuffer_sbuf_p1_rdat_1496};
  assign _zz_shareBuffer_sbuf_p1_rdat_1605 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1606 = {_zz_shareBuffer_sbuf_p1_rdat_1607,_zz_shareBuffer_sbuf_p1_rdat_1608};
  assign _zz_shareBuffer_sbuf_p1_rdat_1715 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1716 = {_zz_shareBuffer_sbuf_p1_rdat_1717,_zz_shareBuffer_sbuf_p1_rdat_1718};
  assign _zz_shareBuffer_sbuf_p1_rdat_32 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_33 = {_zz_shareBuffer_sbuf_p1_rdat_34,_zz_shareBuffer_sbuf_p1_rdat_35};
  assign _zz_shareBuffer_sbuf_p1_rdat_141 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_142 = {_zz_shareBuffer_sbuf_p1_rdat_143,_zz_shareBuffer_sbuf_p1_rdat_144};
  assign _zz_shareBuffer_sbuf_p1_rdat_252 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_253 = {_zz_shareBuffer_sbuf_p1_rdat_254,_zz_shareBuffer_sbuf_p1_rdat_255};
  assign _zz_shareBuffer_sbuf_p1_rdat_363 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_364 = {_zz_shareBuffer_sbuf_p1_rdat_365,_zz_shareBuffer_sbuf_p1_rdat_366};
  assign _zz_shareBuffer_sbuf_p1_rdat_476 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_477 = {_zz_shareBuffer_sbuf_p1_rdat_478,_zz_shareBuffer_sbuf_p1_rdat_479};
  assign _zz_shareBuffer_sbuf_p1_rdat_589 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_590 = {_zz_shareBuffer_sbuf_p1_rdat_591,_zz_shareBuffer_sbuf_p1_rdat_592};
  assign _zz_shareBuffer_sbuf_p1_rdat_702 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_703 = {_zz_shareBuffer_sbuf_p1_rdat_704,_zz_shareBuffer_sbuf_p1_rdat_705};
  assign _zz_shareBuffer_sbuf_p1_rdat_815 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_816 = {_zz_shareBuffer_sbuf_p1_rdat_817,_zz_shareBuffer_sbuf_p1_rdat_818};
  assign _zz_shareBuffer_sbuf_p1_rdat_930 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_931 = {_zz_shareBuffer_sbuf_p1_rdat_932,_zz_shareBuffer_sbuf_p1_rdat_933};
  assign _zz_shareBuffer_sbuf_p1_rdat_1043 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1044 = {_zz_shareBuffer_sbuf_p1_rdat_1045,_zz_shareBuffer_sbuf_p1_rdat_1046};
  assign _zz_shareBuffer_sbuf_p1_rdat_1157 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1158 = {_zz_shareBuffer_sbuf_p1_rdat_1159,_zz_shareBuffer_sbuf_p1_rdat_1160};
  assign _zz_shareBuffer_sbuf_p1_rdat_1270 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1271 = {_zz_shareBuffer_sbuf_p1_rdat_1272,_zz_shareBuffer_sbuf_p1_rdat_1273};
  assign _zz_shareBuffer_sbuf_p1_rdat_1383 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1384 = {_zz_shareBuffer_sbuf_p1_rdat_1385,_zz_shareBuffer_sbuf_p1_rdat_1386};
  assign _zz_shareBuffer_sbuf_p1_rdat_1495 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1496 = {_zz_shareBuffer_sbuf_p1_rdat_1497,_zz_shareBuffer_sbuf_p1_rdat_1498};
  assign _zz_shareBuffer_sbuf_p1_rdat_1607 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1608 = {_zz_shareBuffer_sbuf_p1_rdat_1609,_zz_shareBuffer_sbuf_p1_rdat_1610};
  assign _zz_shareBuffer_sbuf_p1_rdat_1717 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1718 = {_zz_shareBuffer_sbuf_p1_rdat_1719,_zz_shareBuffer_sbuf_p1_rdat_1720};
  assign _zz_shareBuffer_sbuf_p1_rdat_34 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_35 = {_zz_shareBuffer_sbuf_p1_rdat_36,_zz_shareBuffer_sbuf_p1_rdat_37};
  assign _zz_shareBuffer_sbuf_p1_rdat_143 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_144 = {_zz_shareBuffer_sbuf_p1_rdat_145,_zz_shareBuffer_sbuf_p1_rdat_146};
  assign _zz_shareBuffer_sbuf_p1_rdat_254 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_255 = {_zz_shareBuffer_sbuf_p1_rdat_256,_zz_shareBuffer_sbuf_p1_rdat_257};
  assign _zz_shareBuffer_sbuf_p1_rdat_365 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_366 = {_zz_shareBuffer_sbuf_p1_rdat_367,_zz_shareBuffer_sbuf_p1_rdat_368};
  assign _zz_shareBuffer_sbuf_p1_rdat_478 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_479 = {_zz_shareBuffer_sbuf_p1_rdat_480,_zz_shareBuffer_sbuf_p1_rdat_481};
  assign _zz_shareBuffer_sbuf_p1_rdat_591 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_592 = {_zz_shareBuffer_sbuf_p1_rdat_593,_zz_shareBuffer_sbuf_p1_rdat_594};
  assign _zz_shareBuffer_sbuf_p1_rdat_704 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_705 = {_zz_shareBuffer_sbuf_p1_rdat_706,_zz_shareBuffer_sbuf_p1_rdat_707};
  assign _zz_shareBuffer_sbuf_p1_rdat_817 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_818 = {_zz_shareBuffer_sbuf_p1_rdat_819,_zz_shareBuffer_sbuf_p1_rdat_820};
  assign _zz_shareBuffer_sbuf_p1_rdat_932 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_933 = {_zz_shareBuffer_sbuf_p1_rdat_934,_zz_shareBuffer_sbuf_p1_rdat_935};
  assign _zz_shareBuffer_sbuf_p1_rdat_1045 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1046 = {_zz_shareBuffer_sbuf_p1_rdat_1047,_zz_shareBuffer_sbuf_p1_rdat_1048};
  assign _zz_shareBuffer_sbuf_p1_rdat_1159 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1160 = {_zz_shareBuffer_sbuf_p1_rdat_1161,_zz_shareBuffer_sbuf_p1_rdat_1162};
  assign _zz_shareBuffer_sbuf_p1_rdat_1272 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1273 = {_zz_shareBuffer_sbuf_p1_rdat_1274,_zz_shareBuffer_sbuf_p1_rdat_1275};
  assign _zz_shareBuffer_sbuf_p1_rdat_1385 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1386 = {_zz_shareBuffer_sbuf_p1_rdat_1387,_zz_shareBuffer_sbuf_p1_rdat_1388};
  assign _zz_shareBuffer_sbuf_p1_rdat_1497 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1498 = {_zz_shareBuffer_sbuf_p1_rdat_1499,_zz_shareBuffer_sbuf_p1_rdat_1500};
  assign _zz_shareBuffer_sbuf_p1_rdat_1609 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1610 = {_zz_shareBuffer_sbuf_p1_rdat_1611,_zz_shareBuffer_sbuf_p1_rdat_1612};
  assign _zz_shareBuffer_sbuf_p1_rdat_1719 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1720 = {_zz_shareBuffer_sbuf_p1_rdat_1721,_zz_shareBuffer_sbuf_p1_rdat_1722};
  assign _zz_shareBuffer_sbuf_p1_rdat_36 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_37 = {_zz_shareBuffer_sbuf_p1_rdat_38,_zz_shareBuffer_sbuf_p1_rdat_39};
  assign _zz_shareBuffer_sbuf_p1_rdat_145 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_146 = {_zz_shareBuffer_sbuf_p1_rdat_147,_zz_shareBuffer_sbuf_p1_rdat_148};
  assign _zz_shareBuffer_sbuf_p1_rdat_256 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_257 = {_zz_shareBuffer_sbuf_p1_rdat_258,_zz_shareBuffer_sbuf_p1_rdat_259};
  assign _zz_shareBuffer_sbuf_p1_rdat_367 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_368 = {_zz_shareBuffer_sbuf_p1_rdat_369,_zz_shareBuffer_sbuf_p1_rdat_370};
  assign _zz_shareBuffer_sbuf_p1_rdat_480 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_481 = {_zz_shareBuffer_sbuf_p1_rdat_482,_zz_shareBuffer_sbuf_p1_rdat_483};
  assign _zz_shareBuffer_sbuf_p1_rdat_593 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_594 = {_zz_shareBuffer_sbuf_p1_rdat_595,_zz_shareBuffer_sbuf_p1_rdat_596};
  assign _zz_shareBuffer_sbuf_p1_rdat_706 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_707 = {_zz_shareBuffer_sbuf_p1_rdat_708,_zz_shareBuffer_sbuf_p1_rdat_709};
  assign _zz_shareBuffer_sbuf_p1_rdat_819 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_820 = {_zz_shareBuffer_sbuf_p1_rdat_821,_zz_shareBuffer_sbuf_p1_rdat_822};
  assign _zz_shareBuffer_sbuf_p1_rdat_934 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_935 = {_zz_shareBuffer_sbuf_p1_rdat_936,_zz_shareBuffer_sbuf_p1_rdat_937};
  assign _zz_shareBuffer_sbuf_p1_rdat_1047 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1048 = {_zz_shareBuffer_sbuf_p1_rdat_1049,_zz_shareBuffer_sbuf_p1_rdat_1050};
  assign _zz_shareBuffer_sbuf_p1_rdat_1161 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1162 = {_zz_shareBuffer_sbuf_p1_rdat_1163,_zz_shareBuffer_sbuf_p1_rdat_1164};
  assign _zz_shareBuffer_sbuf_p1_rdat_1274 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1275 = {_zz_shareBuffer_sbuf_p1_rdat_1276,_zz_shareBuffer_sbuf_p1_rdat_1277};
  assign _zz_shareBuffer_sbuf_p1_rdat_1387 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1388 = {_zz_shareBuffer_sbuf_p1_rdat_1389,_zz_shareBuffer_sbuf_p1_rdat_1390};
  assign _zz_shareBuffer_sbuf_p1_rdat_1499 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1500 = {_zz_shareBuffer_sbuf_p1_rdat_1501,_zz_shareBuffer_sbuf_p1_rdat_1502};
  assign _zz_shareBuffer_sbuf_p1_rdat_1611 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1612 = {_zz_shareBuffer_sbuf_p1_rdat_1613,_zz_shareBuffer_sbuf_p1_rdat_1614};
  assign _zz_shareBuffer_sbuf_p1_rdat_1721 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1722 = {_zz_shareBuffer_sbuf_p1_rdat_1723,_zz_shareBuffer_sbuf_p1_rdat_1724};
  assign _zz_shareBuffer_sbuf_p1_rdat_38 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_39 = {_zz_shareBuffer_sbuf_p1_rdat_40,_zz_shareBuffer_sbuf_p1_rdat_41};
  assign _zz_shareBuffer_sbuf_p1_rdat_147 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_148 = {_zz_shareBuffer_sbuf_p1_rdat_149,_zz_shareBuffer_sbuf_p1_rdat_150};
  assign _zz_shareBuffer_sbuf_p1_rdat_258 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_259 = {_zz_shareBuffer_sbuf_p1_rdat_260,_zz_shareBuffer_sbuf_p1_rdat_261};
  assign _zz_shareBuffer_sbuf_p1_rdat_369 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_370 = {_zz_shareBuffer_sbuf_p1_rdat_371,_zz_shareBuffer_sbuf_p1_rdat_372};
  assign _zz_shareBuffer_sbuf_p1_rdat_482 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_483 = {_zz_shareBuffer_sbuf_p1_rdat_484,_zz_shareBuffer_sbuf_p1_rdat_485};
  assign _zz_shareBuffer_sbuf_p1_rdat_595 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_596 = {_zz_shareBuffer_sbuf_p1_rdat_597,_zz_shareBuffer_sbuf_p1_rdat_598};
  assign _zz_shareBuffer_sbuf_p1_rdat_708 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_709 = {_zz_shareBuffer_sbuf_p1_rdat_710,_zz_shareBuffer_sbuf_p1_rdat_711};
  assign _zz_shareBuffer_sbuf_p1_rdat_821 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_822 = {_zz_shareBuffer_sbuf_p1_rdat_823,_zz_shareBuffer_sbuf_p1_rdat_824};
  assign _zz_shareBuffer_sbuf_p1_rdat_936 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_937 = {_zz_shareBuffer_sbuf_p1_rdat_938,_zz_shareBuffer_sbuf_p1_rdat_939};
  assign _zz_shareBuffer_sbuf_p1_rdat_1049 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1050 = {_zz_shareBuffer_sbuf_p1_rdat_1051,_zz_shareBuffer_sbuf_p1_rdat_1052};
  assign _zz_shareBuffer_sbuf_p1_rdat_1163 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1164 = {_zz_shareBuffer_sbuf_p1_rdat_1165,_zz_shareBuffer_sbuf_p1_rdat_1166};
  assign _zz_shareBuffer_sbuf_p1_rdat_1276 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1277 = {_zz_shareBuffer_sbuf_p1_rdat_1278,_zz_shareBuffer_sbuf_p1_rdat_1279};
  assign _zz_shareBuffer_sbuf_p1_rdat_1389 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1390 = {_zz_shareBuffer_sbuf_p1_rdat_1391,_zz_shareBuffer_sbuf_p1_rdat_1392};
  assign _zz_shareBuffer_sbuf_p1_rdat_1501 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1502 = {_zz_shareBuffer_sbuf_p1_rdat_1503,_zz_shareBuffer_sbuf_p1_rdat_1504};
  assign _zz_shareBuffer_sbuf_p1_rdat_1613 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1614 = {_zz_shareBuffer_sbuf_p1_rdat_1615,_zz_shareBuffer_sbuf_p1_rdat_1616};
  assign _zz_shareBuffer_sbuf_p1_rdat_1723 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1724 = {_zz_shareBuffer_sbuf_p1_rdat_1725,_zz_shareBuffer_sbuf_p1_rdat_1726};
  assign _zz_shareBuffer_sbuf_p1_rdat_40 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_41 = {_zz_shareBuffer_sbuf_p1_rdat_42,_zz_shareBuffer_sbuf_p1_rdat_43};
  assign _zz_shareBuffer_sbuf_p1_rdat_149 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_150 = {_zz_shareBuffer_sbuf_p1_rdat_151,_zz_shareBuffer_sbuf_p1_rdat_152};
  assign _zz_shareBuffer_sbuf_p1_rdat_260 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_261 = {_zz_shareBuffer_sbuf_p1_rdat_262,_zz_shareBuffer_sbuf_p1_rdat_263};
  assign _zz_shareBuffer_sbuf_p1_rdat_371 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_372 = {_zz_shareBuffer_sbuf_p1_rdat_373,_zz_shareBuffer_sbuf_p1_rdat_374};
  assign _zz_shareBuffer_sbuf_p1_rdat_484 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_485 = {_zz_shareBuffer_sbuf_p1_rdat_486,_zz_shareBuffer_sbuf_p1_rdat_487};
  assign _zz_shareBuffer_sbuf_p1_rdat_597 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_598 = {_zz_shareBuffer_sbuf_p1_rdat_599,_zz_shareBuffer_sbuf_p1_rdat_600};
  assign _zz_shareBuffer_sbuf_p1_rdat_710 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_711 = {_zz_shareBuffer_sbuf_p1_rdat_712,_zz_shareBuffer_sbuf_p1_rdat_713};
  assign _zz_shareBuffer_sbuf_p1_rdat_823 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_824 = {_zz_shareBuffer_sbuf_p1_rdat_825,_zz_shareBuffer_sbuf_p1_rdat_826};
  assign _zz_shareBuffer_sbuf_p1_rdat_938 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_939 = {_zz_shareBuffer_sbuf_p1_rdat_940,_zz_shareBuffer_sbuf_p1_rdat_941};
  assign _zz_shareBuffer_sbuf_p1_rdat_1051 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1052 = {_zz_shareBuffer_sbuf_p1_rdat_1053,_zz_shareBuffer_sbuf_p1_rdat_1054};
  assign _zz_shareBuffer_sbuf_p1_rdat_1165 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1166 = {_zz_shareBuffer_sbuf_p1_rdat_1167,_zz_shareBuffer_sbuf_p1_rdat_1168};
  assign _zz_shareBuffer_sbuf_p1_rdat_1278 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1279 = {_zz_shareBuffer_sbuf_p1_rdat_1280,_zz_shareBuffer_sbuf_p1_rdat_1281};
  assign _zz_shareBuffer_sbuf_p1_rdat_1391 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1392 = {_zz_shareBuffer_sbuf_p1_rdat_1393,_zz_shareBuffer_sbuf_p1_rdat_1394};
  assign _zz_shareBuffer_sbuf_p1_rdat_1503 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1504 = {_zz_shareBuffer_sbuf_p1_rdat_1505,_zz_shareBuffer_sbuf_p1_rdat_1506};
  assign _zz_shareBuffer_sbuf_p1_rdat_1615 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1616 = {_zz_shareBuffer_sbuf_p1_rdat_1617,_zz_shareBuffer_sbuf_p1_rdat_1618};
  assign _zz_shareBuffer_sbuf_p1_rdat_1725 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1726 = {_zz_shareBuffer_sbuf_p1_rdat_1727,_zz_shareBuffer_sbuf_p1_rdat_1728};
  assign _zz_shareBuffer_sbuf_p1_rdat_42 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_43 = {_zz_shareBuffer_sbuf_p1_rdat_44,_zz_shareBuffer_sbuf_p1_rdat_45};
  assign _zz_shareBuffer_sbuf_p1_rdat_151 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_152 = {_zz_shareBuffer_sbuf_p1_rdat_153,_zz_shareBuffer_sbuf_p1_rdat_154};
  assign _zz_shareBuffer_sbuf_p1_rdat_262 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_263 = {_zz_shareBuffer_sbuf_p1_rdat_264,_zz_shareBuffer_sbuf_p1_rdat_265};
  assign _zz_shareBuffer_sbuf_p1_rdat_373 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_374 = {_zz_shareBuffer_sbuf_p1_rdat_375,_zz_shareBuffer_sbuf_p1_rdat_376};
  assign _zz_shareBuffer_sbuf_p1_rdat_486 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_487 = {_zz_shareBuffer_sbuf_p1_rdat_488,_zz_shareBuffer_sbuf_p1_rdat_489};
  assign _zz_shareBuffer_sbuf_p1_rdat_599 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_600 = {_zz_shareBuffer_sbuf_p1_rdat_601,_zz_shareBuffer_sbuf_p1_rdat_602};
  assign _zz_shareBuffer_sbuf_p1_rdat_712 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_713 = {_zz_shareBuffer_sbuf_p1_rdat_714,_zz_shareBuffer_sbuf_p1_rdat_715};
  assign _zz_shareBuffer_sbuf_p1_rdat_825 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_826 = {_zz_shareBuffer_sbuf_p1_rdat_827,_zz_shareBuffer_sbuf_p1_rdat_828};
  assign _zz_shareBuffer_sbuf_p1_rdat_940 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_941 = {_zz_shareBuffer_sbuf_p1_rdat_942,_zz_shareBuffer_sbuf_p1_rdat_943};
  assign _zz_shareBuffer_sbuf_p1_rdat_1053 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1054 = {_zz_shareBuffer_sbuf_p1_rdat_1055,_zz_shareBuffer_sbuf_p1_rdat_1056};
  assign _zz_shareBuffer_sbuf_p1_rdat_1167 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1168 = {_zz_shareBuffer_sbuf_p1_rdat_1169,_zz_shareBuffer_sbuf_p1_rdat_1170};
  assign _zz_shareBuffer_sbuf_p1_rdat_1280 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1281 = {_zz_shareBuffer_sbuf_p1_rdat_1282,_zz_shareBuffer_sbuf_p1_rdat_1283};
  assign _zz_shareBuffer_sbuf_p1_rdat_1393 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1394 = {_zz_shareBuffer_sbuf_p1_rdat_1395,_zz_shareBuffer_sbuf_p1_rdat_1396};
  assign _zz_shareBuffer_sbuf_p1_rdat_1505 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1506 = {_zz_shareBuffer_sbuf_p1_rdat_1507,_zz_shareBuffer_sbuf_p1_rdat_1508};
  assign _zz_shareBuffer_sbuf_p1_rdat_1617 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1618 = {_zz_shareBuffer_sbuf_p1_rdat_1619,_zz_shareBuffer_sbuf_p1_rdat_1620};
  assign _zz_shareBuffer_sbuf_p1_rdat_1727 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1728 = {_zz_shareBuffer_sbuf_p1_rdat_1729,_zz_shareBuffer_sbuf_p1_rdat_1730};
  assign _zz_shareBuffer_sbuf_p1_rdat_44 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_45 = {_zz_shareBuffer_sbuf_p1_rdat_46,_zz_shareBuffer_sbuf_p1_rdat_47};
  assign _zz_shareBuffer_sbuf_p1_rdat_153 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_154 = {_zz_shareBuffer_sbuf_p1_rdat_155,_zz_shareBuffer_sbuf_p1_rdat_156};
  assign _zz_shareBuffer_sbuf_p1_rdat_264 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_265 = {_zz_shareBuffer_sbuf_p1_rdat_266,_zz_shareBuffer_sbuf_p1_rdat_267};
  assign _zz_shareBuffer_sbuf_p1_rdat_375 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_376 = {_zz_shareBuffer_sbuf_p1_rdat_377,_zz_shareBuffer_sbuf_p1_rdat_378};
  assign _zz_shareBuffer_sbuf_p1_rdat_488 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_489 = {_zz_shareBuffer_sbuf_p1_rdat_490,_zz_shareBuffer_sbuf_p1_rdat_491};
  assign _zz_shareBuffer_sbuf_p1_rdat_601 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_602 = {_zz_shareBuffer_sbuf_p1_rdat_603,_zz_shareBuffer_sbuf_p1_rdat_604};
  assign _zz_shareBuffer_sbuf_p1_rdat_714 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_715 = {_zz_shareBuffer_sbuf_p1_rdat_716,_zz_shareBuffer_sbuf_p1_rdat_717};
  assign _zz_shareBuffer_sbuf_p1_rdat_827 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_828 = {_zz_shareBuffer_sbuf_p1_rdat_829,_zz_shareBuffer_sbuf_p1_rdat_830};
  assign _zz_shareBuffer_sbuf_p1_rdat_942 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_943 = {_zz_shareBuffer_sbuf_p1_rdat_944,_zz_shareBuffer_sbuf_p1_rdat_945};
  assign _zz_shareBuffer_sbuf_p1_rdat_1055 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1056 = {_zz_shareBuffer_sbuf_p1_rdat_1057,_zz_shareBuffer_sbuf_p1_rdat_1058};
  assign _zz_shareBuffer_sbuf_p1_rdat_1169 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1170 = {_zz_shareBuffer_sbuf_p1_rdat_1171,_zz_shareBuffer_sbuf_p1_rdat_1172};
  assign _zz_shareBuffer_sbuf_p1_rdat_1282 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1283 = {_zz_shareBuffer_sbuf_p1_rdat_1284,_zz_shareBuffer_sbuf_p1_rdat_1285};
  assign _zz_shareBuffer_sbuf_p1_rdat_1395 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1396 = {_zz_shareBuffer_sbuf_p1_rdat_1397,_zz_shareBuffer_sbuf_p1_rdat_1398};
  assign _zz_shareBuffer_sbuf_p1_rdat_1507 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1508 = {_zz_shareBuffer_sbuf_p1_rdat_1509,_zz_shareBuffer_sbuf_p1_rdat_1510};
  assign _zz_shareBuffer_sbuf_p1_rdat_1619 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1620 = {_zz_shareBuffer_sbuf_p1_rdat_1621,_zz_shareBuffer_sbuf_p1_rdat_1622};
  assign _zz_shareBuffer_sbuf_p1_rdat_1729 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1730 = {_zz_shareBuffer_sbuf_p1_rdat_1731,_zz_shareBuffer_sbuf_p1_rdat_1732};
  assign _zz_shareBuffer_sbuf_p1_rdat_46 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_47 = {_zz_shareBuffer_sbuf_p1_rdat_48,_zz_shareBuffer_sbuf_p1_rdat_49};
  assign _zz_shareBuffer_sbuf_p1_rdat_155 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_156 = {_zz_shareBuffer_sbuf_p1_rdat_157,_zz_shareBuffer_sbuf_p1_rdat_158};
  assign _zz_shareBuffer_sbuf_p1_rdat_266 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_267 = {_zz_shareBuffer_sbuf_p1_rdat_268,_zz_shareBuffer_sbuf_p1_rdat_269};
  assign _zz_shareBuffer_sbuf_p1_rdat_377 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_378 = {_zz_shareBuffer_sbuf_p1_rdat_379,_zz_shareBuffer_sbuf_p1_rdat_380};
  assign _zz_shareBuffer_sbuf_p1_rdat_490 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_491 = {_zz_shareBuffer_sbuf_p1_rdat_492,_zz_shareBuffer_sbuf_p1_rdat_493};
  assign _zz_shareBuffer_sbuf_p1_rdat_603 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_604 = {_zz_shareBuffer_sbuf_p1_rdat_605,_zz_shareBuffer_sbuf_p1_rdat_606};
  assign _zz_shareBuffer_sbuf_p1_rdat_716 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_717 = {_zz_shareBuffer_sbuf_p1_rdat_718,_zz_shareBuffer_sbuf_p1_rdat_719};
  assign _zz_shareBuffer_sbuf_p1_rdat_829 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_830 = {_zz_shareBuffer_sbuf_p1_rdat_831,_zz_shareBuffer_sbuf_p1_rdat_832};
  assign _zz_shareBuffer_sbuf_p1_rdat_944 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_945 = {_zz_shareBuffer_sbuf_p1_rdat_946,_zz_shareBuffer_sbuf_p1_rdat_947};
  assign _zz_shareBuffer_sbuf_p1_rdat_1057 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1058 = {_zz_shareBuffer_sbuf_p1_rdat_1059,_zz_shareBuffer_sbuf_p1_rdat_1060};
  assign _zz_shareBuffer_sbuf_p1_rdat_1171 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1172 = {_zz_shareBuffer_sbuf_p1_rdat_1173,_zz_shareBuffer_sbuf_p1_rdat_1174};
  assign _zz_shareBuffer_sbuf_p1_rdat_1284 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1285 = {_zz_shareBuffer_sbuf_p1_rdat_1286,_zz_shareBuffer_sbuf_p1_rdat_1287};
  assign _zz_shareBuffer_sbuf_p1_rdat_1397 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1398 = {_zz_shareBuffer_sbuf_p1_rdat_1399,_zz_shareBuffer_sbuf_p1_rdat_1400};
  assign _zz_shareBuffer_sbuf_p1_rdat_1509 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1510 = {_zz_shareBuffer_sbuf_p1_rdat_1511,_zz_shareBuffer_sbuf_p1_rdat_1512};
  assign _zz_shareBuffer_sbuf_p1_rdat_1621 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1622 = {_zz_shareBuffer_sbuf_p1_rdat_1623,_zz_shareBuffer_sbuf_p1_rdat_1624};
  assign _zz_shareBuffer_sbuf_p1_rdat_1731 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1732 = {_zz_shareBuffer_sbuf_p1_rdat_1733,_zz_shareBuffer_sbuf_p1_rdat_1734};
  assign _zz_shareBuffer_sbuf_p1_rdat_48 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_49 = {_zz_shareBuffer_sbuf_p1_rdat_50,_zz_shareBuffer_sbuf_p1_rdat_51};
  assign _zz_shareBuffer_sbuf_p1_rdat_157 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_158 = {_zz_shareBuffer_sbuf_p1_rdat_159,_zz_shareBuffer_sbuf_p1_rdat_160};
  assign _zz_shareBuffer_sbuf_p1_rdat_268 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_269 = {_zz_shareBuffer_sbuf_p1_rdat_270,_zz_shareBuffer_sbuf_p1_rdat_271};
  assign _zz_shareBuffer_sbuf_p1_rdat_379 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_380 = {_zz_shareBuffer_sbuf_p1_rdat_381,_zz_shareBuffer_sbuf_p1_rdat_382};
  assign _zz_shareBuffer_sbuf_p1_rdat_492 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_493 = {_zz_shareBuffer_sbuf_p1_rdat_494,_zz_shareBuffer_sbuf_p1_rdat_495};
  assign _zz_shareBuffer_sbuf_p1_rdat_605 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_606 = {_zz_shareBuffer_sbuf_p1_rdat_607,_zz_shareBuffer_sbuf_p1_rdat_608};
  assign _zz_shareBuffer_sbuf_p1_rdat_718 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_719 = {_zz_shareBuffer_sbuf_p1_rdat_720,_zz_shareBuffer_sbuf_p1_rdat_721};
  assign _zz_shareBuffer_sbuf_p1_rdat_831 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_832 = {_zz_shareBuffer_sbuf_p1_rdat_833,_zz_shareBuffer_sbuf_p1_rdat_834};
  assign _zz_shareBuffer_sbuf_p1_rdat_946 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_947 = {_zz_shareBuffer_sbuf_p1_rdat_948,_zz_shareBuffer_sbuf_p1_rdat_949};
  assign _zz_shareBuffer_sbuf_p1_rdat_1059 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1060 = {_zz_shareBuffer_sbuf_p1_rdat_1061,_zz_shareBuffer_sbuf_p1_rdat_1062};
  assign _zz_shareBuffer_sbuf_p1_rdat_1173 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1174 = {_zz_shareBuffer_sbuf_p1_rdat_1175,_zz_shareBuffer_sbuf_p1_rdat_1176};
  assign _zz_shareBuffer_sbuf_p1_rdat_1286 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1287 = {_zz_shareBuffer_sbuf_p1_rdat_1288,_zz_shareBuffer_sbuf_p1_rdat_1289};
  assign _zz_shareBuffer_sbuf_p1_rdat_1399 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1400 = {_zz_shareBuffer_sbuf_p1_rdat_1401,_zz_shareBuffer_sbuf_p1_rdat_1402};
  assign _zz_shareBuffer_sbuf_p1_rdat_1511 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1512 = {_zz_shareBuffer_sbuf_p1_rdat_1513,_zz_shareBuffer_sbuf_p1_rdat_1514};
  assign _zz_shareBuffer_sbuf_p1_rdat_1623 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1624 = {_zz_shareBuffer_sbuf_p1_rdat_1625,_zz_shareBuffer_sbuf_p1_rdat_1626};
  assign _zz_shareBuffer_sbuf_p1_rdat_1733 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1734 = {_zz_shareBuffer_sbuf_p1_rdat_1735,_zz_shareBuffer_sbuf_p1_rdat_1736};
  assign _zz_shareBuffer_sbuf_p1_rdat_50 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_51 = {_zz_shareBuffer_sbuf_p1_rdat_52,_zz_shareBuffer_sbuf_p1_rdat_53};
  assign _zz_shareBuffer_sbuf_p1_rdat_159 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_160 = {_zz_shareBuffer_sbuf_p1_rdat_161,_zz_shareBuffer_sbuf_p1_rdat_162};
  assign _zz_shareBuffer_sbuf_p1_rdat_270 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_271 = {_zz_shareBuffer_sbuf_p1_rdat_272,_zz_shareBuffer_sbuf_p1_rdat_273};
  assign _zz_shareBuffer_sbuf_p1_rdat_381 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_382 = {_zz_shareBuffer_sbuf_p1_rdat_383,_zz_shareBuffer_sbuf_p1_rdat_384};
  assign _zz_shareBuffer_sbuf_p1_rdat_494 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_495 = {_zz_shareBuffer_sbuf_p1_rdat_496,_zz_shareBuffer_sbuf_p1_rdat_497};
  assign _zz_shareBuffer_sbuf_p1_rdat_607 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_608 = {_zz_shareBuffer_sbuf_p1_rdat_609,_zz_shareBuffer_sbuf_p1_rdat_610};
  assign _zz_shareBuffer_sbuf_p1_rdat_720 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_721 = {_zz_shareBuffer_sbuf_p1_rdat_722,_zz_shareBuffer_sbuf_p1_rdat_723};
  assign _zz_shareBuffer_sbuf_p1_rdat_833 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_834 = {_zz_shareBuffer_sbuf_p1_rdat_835,_zz_shareBuffer_sbuf_p1_rdat_836};
  assign _zz_shareBuffer_sbuf_p1_rdat_948 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_949 = {_zz_shareBuffer_sbuf_p1_rdat_950,_zz_shareBuffer_sbuf_p1_rdat_951};
  assign _zz_shareBuffer_sbuf_p1_rdat_1061 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1062 = {_zz_shareBuffer_sbuf_p1_rdat_1063,_zz_shareBuffer_sbuf_p1_rdat_1064};
  assign _zz_shareBuffer_sbuf_p1_rdat_1175 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1176 = {_zz_shareBuffer_sbuf_p1_rdat_1177,_zz_shareBuffer_sbuf_p1_rdat_1178};
  assign _zz_shareBuffer_sbuf_p1_rdat_1288 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1289 = {_zz_shareBuffer_sbuf_p1_rdat_1290,_zz_shareBuffer_sbuf_p1_rdat_1291};
  assign _zz_shareBuffer_sbuf_p1_rdat_1401 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1402 = {_zz_shareBuffer_sbuf_p1_rdat_1403,_zz_shareBuffer_sbuf_p1_rdat_1404};
  assign _zz_shareBuffer_sbuf_p1_rdat_1513 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1514 = {_zz_shareBuffer_sbuf_p1_rdat_1515,_zz_shareBuffer_sbuf_p1_rdat_1516};
  assign _zz_shareBuffer_sbuf_p1_rdat_1625 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1626 = {_zz_shareBuffer_sbuf_p1_rdat_1627,_zz_shareBuffer_sbuf_p1_rdat_1628};
  assign _zz_shareBuffer_sbuf_p1_rdat_1735 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1736 = {_zz_shareBuffer_sbuf_p1_rdat_1737,_zz_shareBuffer_sbuf_p1_rdat_1738};
  assign _zz_shareBuffer_sbuf_p1_rdat_52 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_53 = {_zz_shareBuffer_sbuf_p1_rdat_54,_zz_shareBuffer_sbuf_p1_rdat_55};
  assign _zz_shareBuffer_sbuf_p1_rdat_161 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_162 = {_zz_shareBuffer_sbuf_p1_rdat_163,_zz_shareBuffer_sbuf_p1_rdat_164};
  assign _zz_shareBuffer_sbuf_p1_rdat_272 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_273 = {_zz_shareBuffer_sbuf_p1_rdat_274,_zz_shareBuffer_sbuf_p1_rdat_275};
  assign _zz_shareBuffer_sbuf_p1_rdat_383 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_384 = {_zz_shareBuffer_sbuf_p1_rdat_385,_zz_shareBuffer_sbuf_p1_rdat_386};
  assign _zz_shareBuffer_sbuf_p1_rdat_496 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_497 = {_zz_shareBuffer_sbuf_p1_rdat_498,_zz_shareBuffer_sbuf_p1_rdat_499};
  assign _zz_shareBuffer_sbuf_p1_rdat_609 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_610 = {_zz_shareBuffer_sbuf_p1_rdat_611,_zz_shareBuffer_sbuf_p1_rdat_612};
  assign _zz_shareBuffer_sbuf_p1_rdat_722 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_723 = {_zz_shareBuffer_sbuf_p1_rdat_724,_zz_shareBuffer_sbuf_p1_rdat_725};
  assign _zz_shareBuffer_sbuf_p1_rdat_835 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_836 = {_zz_shareBuffer_sbuf_p1_rdat_837,_zz_shareBuffer_sbuf_p1_rdat_838};
  assign _zz_shareBuffer_sbuf_p1_rdat_950 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_951 = {_zz_shareBuffer_sbuf_p1_rdat_952,_zz_shareBuffer_sbuf_p1_rdat_953};
  assign _zz_shareBuffer_sbuf_p1_rdat_1063 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1064 = {_zz_shareBuffer_sbuf_p1_rdat_1065,_zz_shareBuffer_sbuf_p1_rdat_1066};
  assign _zz_shareBuffer_sbuf_p1_rdat_1177 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1178 = {_zz_shareBuffer_sbuf_p1_rdat_1179,_zz_shareBuffer_sbuf_p1_rdat_1180};
  assign _zz_shareBuffer_sbuf_p1_rdat_1290 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1291 = {_zz_shareBuffer_sbuf_p1_rdat_1292,_zz_shareBuffer_sbuf_p1_rdat_1293};
  assign _zz_shareBuffer_sbuf_p1_rdat_1403 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1404 = {_zz_shareBuffer_sbuf_p1_rdat_1405,_zz_shareBuffer_sbuf_p1_rdat_1406};
  assign _zz_shareBuffer_sbuf_p1_rdat_1515 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1516 = {_zz_shareBuffer_sbuf_p1_rdat_1517,_zz_shareBuffer_sbuf_p1_rdat_1518};
  assign _zz_shareBuffer_sbuf_p1_rdat_1627 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1628 = {_zz_shareBuffer_sbuf_p1_rdat_1629,_zz_shareBuffer_sbuf_p1_rdat_1630};
  assign _zz_shareBuffer_sbuf_p1_rdat_1737 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1738 = {_zz_shareBuffer_sbuf_p1_rdat_1739,_zz_shareBuffer_sbuf_p1_rdat_1740};
  assign _zz_shareBuffer_sbuf_p1_rdat_54 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_55 = {_zz_shareBuffer_sbuf_p1_rdat_56,_zz_shareBuffer_sbuf_p1_rdat_57};
  assign _zz_shareBuffer_sbuf_p1_rdat_163 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_164 = {_zz_shareBuffer_sbuf_p1_rdat_165,_zz_shareBuffer_sbuf_p1_rdat_166};
  assign _zz_shareBuffer_sbuf_p1_rdat_274 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_275 = {_zz_shareBuffer_sbuf_p1_rdat_276,_zz_shareBuffer_sbuf_p1_rdat_277};
  assign _zz_shareBuffer_sbuf_p1_rdat_385 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_386 = {_zz_shareBuffer_sbuf_p1_rdat_387,_zz_shareBuffer_sbuf_p1_rdat_388};
  assign _zz_shareBuffer_sbuf_p1_rdat_498 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_499 = {_zz_shareBuffer_sbuf_p1_rdat_500,_zz_shareBuffer_sbuf_p1_rdat_501};
  assign _zz_shareBuffer_sbuf_p1_rdat_611 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_612 = {_zz_shareBuffer_sbuf_p1_rdat_613,_zz_shareBuffer_sbuf_p1_rdat_614};
  assign _zz_shareBuffer_sbuf_p1_rdat_724 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_725 = {_zz_shareBuffer_sbuf_p1_rdat_726,_zz_shareBuffer_sbuf_p1_rdat_727};
  assign _zz_shareBuffer_sbuf_p1_rdat_837 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_838 = {_zz_shareBuffer_sbuf_p1_rdat_839,_zz_shareBuffer_sbuf_p1_rdat_840};
  assign _zz_shareBuffer_sbuf_p1_rdat_952 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_953 = {_zz_shareBuffer_sbuf_p1_rdat_954,_zz_shareBuffer_sbuf_p1_rdat_955};
  assign _zz_shareBuffer_sbuf_p1_rdat_1065 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1066 = {_zz_shareBuffer_sbuf_p1_rdat_1067,_zz_shareBuffer_sbuf_p1_rdat_1068};
  assign _zz_shareBuffer_sbuf_p1_rdat_1179 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1180 = {_zz_shareBuffer_sbuf_p1_rdat_1181,_zz_shareBuffer_sbuf_p1_rdat_1182};
  assign _zz_shareBuffer_sbuf_p1_rdat_1292 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1293 = {_zz_shareBuffer_sbuf_p1_rdat_1294,_zz_shareBuffer_sbuf_p1_rdat_1295};
  assign _zz_shareBuffer_sbuf_p1_rdat_1405 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1406 = {_zz_shareBuffer_sbuf_p1_rdat_1407,_zz_shareBuffer_sbuf_p1_rdat_1408};
  assign _zz_shareBuffer_sbuf_p1_rdat_1517 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1518 = {_zz_shareBuffer_sbuf_p1_rdat_1519,_zz_shareBuffer_sbuf_p1_rdat_1520};
  assign _zz_shareBuffer_sbuf_p1_rdat_1629 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1630 = {_zz_shareBuffer_sbuf_p1_rdat_1631,_zz_shareBuffer_sbuf_p1_rdat_1632};
  assign _zz_shareBuffer_sbuf_p1_rdat_1739 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1740 = {_zz_shareBuffer_sbuf_p1_rdat_1741,_zz_shareBuffer_sbuf_p1_rdat_1742};
  assign _zz_shareBuffer_sbuf_p1_rdat_56 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_57 = {_zz_shareBuffer_sbuf_p1_rdat_58,_zz_shareBuffer_sbuf_p1_rdat_59};
  assign _zz_shareBuffer_sbuf_p1_rdat_165 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_166 = {_zz_shareBuffer_sbuf_p1_rdat_167,_zz_shareBuffer_sbuf_p1_rdat_168};
  assign _zz_shareBuffer_sbuf_p1_rdat_276 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_277 = {_zz_shareBuffer_sbuf_p1_rdat_278,_zz_shareBuffer_sbuf_p1_rdat_279};
  assign _zz_shareBuffer_sbuf_p1_rdat_387 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_388 = {_zz_shareBuffer_sbuf_p1_rdat_389,_zz_shareBuffer_sbuf_p1_rdat_390};
  assign _zz_shareBuffer_sbuf_p1_rdat_500 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_501 = {_zz_shareBuffer_sbuf_p1_rdat_502,_zz_shareBuffer_sbuf_p1_rdat_503};
  assign _zz_shareBuffer_sbuf_p1_rdat_613 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_614 = {_zz_shareBuffer_sbuf_p1_rdat_615,_zz_shareBuffer_sbuf_p1_rdat_616};
  assign _zz_shareBuffer_sbuf_p1_rdat_726 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_727 = {_zz_shareBuffer_sbuf_p1_rdat_728,_zz_shareBuffer_sbuf_p1_rdat_729};
  assign _zz_shareBuffer_sbuf_p1_rdat_839 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_840 = {_zz_shareBuffer_sbuf_p1_rdat_841,_zz_shareBuffer_sbuf_p1_rdat_842};
  assign _zz_shareBuffer_sbuf_p1_rdat_954 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_955 = {_zz_shareBuffer_sbuf_p1_rdat_956,_zz_shareBuffer_sbuf_p1_rdat_957};
  assign _zz_shareBuffer_sbuf_p1_rdat_1067 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1068 = {_zz_shareBuffer_sbuf_p1_rdat_1069,_zz_shareBuffer_sbuf_p1_rdat_1070};
  assign _zz_shareBuffer_sbuf_p1_rdat_1181 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1182 = {_zz_shareBuffer_sbuf_p1_rdat_1183,_zz_shareBuffer_sbuf_p1_rdat_1184};
  assign _zz_shareBuffer_sbuf_p1_rdat_1294 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1295 = {_zz_shareBuffer_sbuf_p1_rdat_1296,_zz_shareBuffer_sbuf_p1_rdat_1297};
  assign _zz_shareBuffer_sbuf_p1_rdat_1407 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1408 = {_zz_shareBuffer_sbuf_p1_rdat_1409,_zz_shareBuffer_sbuf_p1_rdat_1410};
  assign _zz_shareBuffer_sbuf_p1_rdat_1519 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1520 = {_zz_shareBuffer_sbuf_p1_rdat_1521,_zz_shareBuffer_sbuf_p1_rdat_1522};
  assign _zz_shareBuffer_sbuf_p1_rdat_1631 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1632 = {_zz_shareBuffer_sbuf_p1_rdat_1633,_zz_shareBuffer_sbuf_p1_rdat_1634};
  assign _zz_shareBuffer_sbuf_p1_rdat_1741 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1742 = {_zz_shareBuffer_sbuf_p1_rdat_1743,_zz_shareBuffer_sbuf_p1_rdat_1744};
  assign _zz_shareBuffer_sbuf_p1_rdat_58 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_59 = {_zz_shareBuffer_sbuf_p1_rdat_60,_zz_shareBuffer_sbuf_p1_rdat_61};
  assign _zz_shareBuffer_sbuf_p1_rdat_167 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_168 = {_zz_shareBuffer_sbuf_p1_rdat_169,_zz_shareBuffer_sbuf_p1_rdat_170};
  assign _zz_shareBuffer_sbuf_p1_rdat_278 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_279 = {_zz_shareBuffer_sbuf_p1_rdat_280,_zz_shareBuffer_sbuf_p1_rdat_281};
  assign _zz_shareBuffer_sbuf_p1_rdat_389 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_390 = {_zz_shareBuffer_sbuf_p1_rdat_391,_zz_shareBuffer_sbuf_p1_rdat_392};
  assign _zz_shareBuffer_sbuf_p1_rdat_502 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_503 = {_zz_shareBuffer_sbuf_p1_rdat_504,_zz_shareBuffer_sbuf_p1_rdat_505};
  assign _zz_shareBuffer_sbuf_p1_rdat_615 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_616 = {_zz_shareBuffer_sbuf_p1_rdat_617,_zz_shareBuffer_sbuf_p1_rdat_618};
  assign _zz_shareBuffer_sbuf_p1_rdat_728 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_729 = {_zz_shareBuffer_sbuf_p1_rdat_730,_zz_shareBuffer_sbuf_p1_rdat_731};
  assign _zz_shareBuffer_sbuf_p1_rdat_841 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_842 = {_zz_shareBuffer_sbuf_p1_rdat_843,_zz_shareBuffer_sbuf_p1_rdat_844};
  assign _zz_shareBuffer_sbuf_p1_rdat_956 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_957 = {_zz_shareBuffer_sbuf_p1_rdat_958,_zz_shareBuffer_sbuf_p1_rdat_959};
  assign _zz_shareBuffer_sbuf_p1_rdat_1069 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1070 = {_zz_shareBuffer_sbuf_p1_rdat_1071,_zz_shareBuffer_sbuf_p1_rdat_1072};
  assign _zz_shareBuffer_sbuf_p1_rdat_1183 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1184 = {_zz_shareBuffer_sbuf_p1_rdat_1185,_zz_shareBuffer_sbuf_p1_rdat_1186};
  assign _zz_shareBuffer_sbuf_p1_rdat_1296 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1297 = {_zz_shareBuffer_sbuf_p1_rdat_1298,_zz_shareBuffer_sbuf_p1_rdat_1299};
  assign _zz_shareBuffer_sbuf_p1_rdat_1409 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1410 = {_zz_shareBuffer_sbuf_p1_rdat_1411,_zz_shareBuffer_sbuf_p1_rdat_1412};
  assign _zz_shareBuffer_sbuf_p1_rdat_1521 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1522 = {_zz_shareBuffer_sbuf_p1_rdat_1523,_zz_shareBuffer_sbuf_p1_rdat_1524};
  assign _zz_shareBuffer_sbuf_p1_rdat_1633 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1634 = {_zz_shareBuffer_sbuf_p1_rdat_1635,_zz_shareBuffer_sbuf_p1_rdat_1636};
  assign _zz_shareBuffer_sbuf_p1_rdat_1743 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1744 = {_zz_shareBuffer_sbuf_p1_rdat_1745,_zz_shareBuffer_sbuf_p1_rdat_1746};
  assign _zz_shareBuffer_sbuf_p1_rdat_60 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_61 = {_zz_shareBuffer_sbuf_p1_rdat_62,_zz_shareBuffer_sbuf_p1_rdat_63};
  assign _zz_shareBuffer_sbuf_p1_rdat_169 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_170 = {_zz_shareBuffer_sbuf_p1_rdat_171,_zz_shareBuffer_sbuf_p1_rdat_172};
  assign _zz_shareBuffer_sbuf_p1_rdat_280 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_281 = {_zz_shareBuffer_sbuf_p1_rdat_282,_zz_shareBuffer_sbuf_p1_rdat_283};
  assign _zz_shareBuffer_sbuf_p1_rdat_391 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_392 = {_zz_shareBuffer_sbuf_p1_rdat_393,_zz_shareBuffer_sbuf_p1_rdat_394};
  assign _zz_shareBuffer_sbuf_p1_rdat_504 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_505 = {_zz_shareBuffer_sbuf_p1_rdat_506,_zz_shareBuffer_sbuf_p1_rdat_507};
  assign _zz_shareBuffer_sbuf_p1_rdat_617 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_618 = {_zz_shareBuffer_sbuf_p1_rdat_619,_zz_shareBuffer_sbuf_p1_rdat_620};
  assign _zz_shareBuffer_sbuf_p1_rdat_730 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_731 = {_zz_shareBuffer_sbuf_p1_rdat_732,_zz_shareBuffer_sbuf_p1_rdat_733};
  assign _zz_shareBuffer_sbuf_p1_rdat_843 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_844 = {_zz_shareBuffer_sbuf_p1_rdat_845,_zz_shareBuffer_sbuf_p1_rdat_846};
  assign _zz_shareBuffer_sbuf_p1_rdat_958 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_959 = {_zz_shareBuffer_sbuf_p1_rdat_960,_zz_shareBuffer_sbuf_p1_rdat_961};
  assign _zz_shareBuffer_sbuf_p1_rdat_1071 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1072 = {_zz_shareBuffer_sbuf_p1_rdat_1073,_zz_shareBuffer_sbuf_p1_rdat_1074};
  assign _zz_shareBuffer_sbuf_p1_rdat_1185 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1186 = {_zz_shareBuffer_sbuf_p1_rdat_1187,_zz_shareBuffer_sbuf_p1_rdat_1188};
  assign _zz_shareBuffer_sbuf_p1_rdat_1298 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1299 = {_zz_shareBuffer_sbuf_p1_rdat_1300,_zz_shareBuffer_sbuf_p1_rdat_1301};
  assign _zz_shareBuffer_sbuf_p1_rdat_1411 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1412 = {_zz_shareBuffer_sbuf_p1_rdat_1413,_zz_shareBuffer_sbuf_p1_rdat_1414};
  assign _zz_shareBuffer_sbuf_p1_rdat_1523 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1524 = {_zz_shareBuffer_sbuf_p1_rdat_1525,_zz_shareBuffer_sbuf_p1_rdat_1526};
  assign _zz_shareBuffer_sbuf_p1_rdat_1635 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1636 = {_zz_shareBuffer_sbuf_p1_rdat_1637,_zz_shareBuffer_sbuf_p1_rdat_1638};
  assign _zz_shareBuffer_sbuf_p1_rdat_1745 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1746 = {_zz_shareBuffer_sbuf_p1_rdat_1747,_zz_shareBuffer_sbuf_p1_rdat_1748};
  assign _zz_shareBuffer_sbuf_p1_rdat_62 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_63 = {_zz_shareBuffer_sbuf_p1_rdat_64,_zz_shareBuffer_sbuf_p1_rdat_65};
  assign _zz_shareBuffer_sbuf_p1_rdat_171 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_172 = {_zz_shareBuffer_sbuf_p1_rdat_173,_zz_shareBuffer_sbuf_p1_rdat_174};
  assign _zz_shareBuffer_sbuf_p1_rdat_282 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_283 = {_zz_shareBuffer_sbuf_p1_rdat_284,_zz_shareBuffer_sbuf_p1_rdat_285};
  assign _zz_shareBuffer_sbuf_p1_rdat_393 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_394 = {_zz_shareBuffer_sbuf_p1_rdat_395,_zz_shareBuffer_sbuf_p1_rdat_396};
  assign _zz_shareBuffer_sbuf_p1_rdat_506 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_507 = {_zz_shareBuffer_sbuf_p1_rdat_508,_zz_shareBuffer_sbuf_p1_rdat_509};
  assign _zz_shareBuffer_sbuf_p1_rdat_619 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_620 = {_zz_shareBuffer_sbuf_p1_rdat_621,_zz_shareBuffer_sbuf_p1_rdat_622};
  assign _zz_shareBuffer_sbuf_p1_rdat_732 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_733 = {_zz_shareBuffer_sbuf_p1_rdat_734,_zz_shareBuffer_sbuf_p1_rdat_735};
  assign _zz_shareBuffer_sbuf_p1_rdat_845 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_846 = {_zz_shareBuffer_sbuf_p1_rdat_847,_zz_shareBuffer_sbuf_p1_rdat_848};
  assign _zz_shareBuffer_sbuf_p1_rdat_960 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_961 = {_zz_shareBuffer_sbuf_p1_rdat_962,_zz_shareBuffer_sbuf_p1_rdat_963};
  assign _zz_shareBuffer_sbuf_p1_rdat_1073 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1074 = {_zz_shareBuffer_sbuf_p1_rdat_1075,_zz_shareBuffer_sbuf_p1_rdat_1076};
  assign _zz_shareBuffer_sbuf_p1_rdat_1187 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1188 = {_zz_shareBuffer_sbuf_p1_rdat_1189,_zz_shareBuffer_sbuf_p1_rdat_1190};
  assign _zz_shareBuffer_sbuf_p1_rdat_1300 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1301 = {_zz_shareBuffer_sbuf_p1_rdat_1302,_zz_shareBuffer_sbuf_p1_rdat_1303};
  assign _zz_shareBuffer_sbuf_p1_rdat_1413 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1414 = {_zz_shareBuffer_sbuf_p1_rdat_1415,_zz_shareBuffer_sbuf_p1_rdat_1416};
  assign _zz_shareBuffer_sbuf_p1_rdat_1525 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1526 = {_zz_shareBuffer_sbuf_p1_rdat_1527,_zz_shareBuffer_sbuf_p1_rdat_1528};
  assign _zz_shareBuffer_sbuf_p1_rdat_1637 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1638 = {_zz_shareBuffer_sbuf_p1_rdat_1639,_zz_shareBuffer_sbuf_p1_rdat_1640};
  assign _zz_shareBuffer_sbuf_p1_rdat_1747 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1748 = {_zz_shareBuffer_sbuf_p1_rdat_1749,_zz_shareBuffer_sbuf_p1_rdat_1750};
  assign _zz_shareBuffer_sbuf_p1_rdat_64 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_65 = {_zz_shareBuffer_sbuf_p1_rdat_66,_zz_shareBuffer_sbuf_p1_rdat_67};
  assign _zz_shareBuffer_sbuf_p1_rdat_173 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_174 = {_zz_shareBuffer_sbuf_p1_rdat_175,_zz_shareBuffer_sbuf_p1_rdat_176};
  assign _zz_shareBuffer_sbuf_p1_rdat_284 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_285 = {_zz_shareBuffer_sbuf_p1_rdat_286,_zz_shareBuffer_sbuf_p1_rdat_287};
  assign _zz_shareBuffer_sbuf_p1_rdat_395 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_396 = {_zz_shareBuffer_sbuf_p1_rdat_397,_zz_shareBuffer_sbuf_p1_rdat_398};
  assign _zz_shareBuffer_sbuf_p1_rdat_508 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_509 = {_zz_shareBuffer_sbuf_p1_rdat_510,_zz_shareBuffer_sbuf_p1_rdat_511};
  assign _zz_shareBuffer_sbuf_p1_rdat_621 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_622 = {_zz_shareBuffer_sbuf_p1_rdat_623,_zz_shareBuffer_sbuf_p1_rdat_624};
  assign _zz_shareBuffer_sbuf_p1_rdat_734 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_735 = {_zz_shareBuffer_sbuf_p1_rdat_736,_zz_shareBuffer_sbuf_p1_rdat_737};
  assign _zz_shareBuffer_sbuf_p1_rdat_847 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_848 = {_zz_shareBuffer_sbuf_p1_rdat_849,_zz_shareBuffer_sbuf_p1_rdat_850};
  assign _zz_shareBuffer_sbuf_p1_rdat_962 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_963 = {_zz_shareBuffer_sbuf_p1_rdat_964,_zz_shareBuffer_sbuf_p1_rdat_965};
  assign _zz_shareBuffer_sbuf_p1_rdat_1075 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1076 = {_zz_shareBuffer_sbuf_p1_rdat_1077,_zz_shareBuffer_sbuf_p1_rdat_1078};
  assign _zz_shareBuffer_sbuf_p1_rdat_1189 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1190 = {_zz_shareBuffer_sbuf_p1_rdat_1191,_zz_shareBuffer_sbuf_p1_rdat_1192};
  assign _zz_shareBuffer_sbuf_p1_rdat_1302 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1303 = {_zz_shareBuffer_sbuf_p1_rdat_1304,_zz_shareBuffer_sbuf_p1_rdat_1305};
  assign _zz_shareBuffer_sbuf_p1_rdat_1415 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1416 = {_zz_shareBuffer_sbuf_p1_rdat_1417,_zz_shareBuffer_sbuf_p1_rdat_1418};
  assign _zz_shareBuffer_sbuf_p1_rdat_1527 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1528 = {_zz_shareBuffer_sbuf_p1_rdat_1529,_zz_shareBuffer_sbuf_p1_rdat_1530};
  assign _zz_shareBuffer_sbuf_p1_rdat_1639 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1640 = {_zz_shareBuffer_sbuf_p1_rdat_1641,_zz_shareBuffer_sbuf_p1_rdat_1642};
  assign _zz_shareBuffer_sbuf_p1_rdat_1749 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1750 = {_zz_shareBuffer_sbuf_p1_rdat_1751,_zz_shareBuffer_sbuf_p1_rdat_1752};
  assign _zz_shareBuffer_sbuf_p1_rdat_66 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_67 = {_zz_shareBuffer_sbuf_p1_rdat_68,_zz_shareBuffer_sbuf_p1_rdat_69};
  assign _zz_shareBuffer_sbuf_p1_rdat_175 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_176 = {_zz_shareBuffer_sbuf_p1_rdat_177,_zz_shareBuffer_sbuf_p1_rdat_178};
  assign _zz_shareBuffer_sbuf_p1_rdat_286 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_287 = {_zz_shareBuffer_sbuf_p1_rdat_288,_zz_shareBuffer_sbuf_p1_rdat_289};
  assign _zz_shareBuffer_sbuf_p1_rdat_397 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_398 = {_zz_shareBuffer_sbuf_p1_rdat_399,_zz_shareBuffer_sbuf_p1_rdat_400};
  assign _zz_shareBuffer_sbuf_p1_rdat_510 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_511 = {_zz_shareBuffer_sbuf_p1_rdat_512,_zz_shareBuffer_sbuf_p1_rdat_513};
  assign _zz_shareBuffer_sbuf_p1_rdat_623 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_624 = {_zz_shareBuffer_sbuf_p1_rdat_625,_zz_shareBuffer_sbuf_p1_rdat_626};
  assign _zz_shareBuffer_sbuf_p1_rdat_736 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_737 = {_zz_shareBuffer_sbuf_p1_rdat_738,_zz_shareBuffer_sbuf_p1_rdat_739};
  assign _zz_shareBuffer_sbuf_p1_rdat_849 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_850 = {_zz_shareBuffer_sbuf_p1_rdat_851,_zz_shareBuffer_sbuf_p1_rdat_852};
  assign _zz_shareBuffer_sbuf_p1_rdat_964 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_965 = {_zz_shareBuffer_sbuf_p1_rdat_966,_zz_shareBuffer_sbuf_p1_rdat_967};
  assign _zz_shareBuffer_sbuf_p1_rdat_1077 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1078 = {_zz_shareBuffer_sbuf_p1_rdat_1079,_zz_shareBuffer_sbuf_p1_rdat_1080};
  assign _zz_shareBuffer_sbuf_p1_rdat_1191 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1192 = {_zz_shareBuffer_sbuf_p1_rdat_1193,_zz_shareBuffer_sbuf_p1_rdat_1194};
  assign _zz_shareBuffer_sbuf_p1_rdat_1304 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1305 = {_zz_shareBuffer_sbuf_p1_rdat_1306,_zz_shareBuffer_sbuf_p1_rdat_1307};
  assign _zz_shareBuffer_sbuf_p1_rdat_1417 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1418 = {_zz_shareBuffer_sbuf_p1_rdat_1419,_zz_shareBuffer_sbuf_p1_rdat_1420};
  assign _zz_shareBuffer_sbuf_p1_rdat_1529 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1530 = {_zz_shareBuffer_sbuf_p1_rdat_1531,_zz_shareBuffer_sbuf_p1_rdat_1532};
  assign _zz_shareBuffer_sbuf_p1_rdat_1641 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1642 = {_zz_shareBuffer_sbuf_p1_rdat_1643,_zz_shareBuffer_sbuf_p1_rdat_1644};
  assign _zz_shareBuffer_sbuf_p1_rdat_1751 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1752 = {_zz_shareBuffer_sbuf_p1_rdat_1753,_zz_shareBuffer_sbuf_p1_rdat_1754};
  assign _zz_shareBuffer_sbuf_p1_rdat_68 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_69 = {_zz_shareBuffer_sbuf_p1_rdat_70,_zz_shareBuffer_sbuf_p1_rdat_71};
  assign _zz_shareBuffer_sbuf_p1_rdat_177 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_178 = {_zz_shareBuffer_sbuf_p1_rdat_179,_zz_shareBuffer_sbuf_p1_rdat_180};
  assign _zz_shareBuffer_sbuf_p1_rdat_288 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_289 = {_zz_shareBuffer_sbuf_p1_rdat_290,_zz_shareBuffer_sbuf_p1_rdat_291};
  assign _zz_shareBuffer_sbuf_p1_rdat_399 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_400 = {_zz_shareBuffer_sbuf_p1_rdat_401,_zz_shareBuffer_sbuf_p1_rdat_402};
  assign _zz_shareBuffer_sbuf_p1_rdat_512 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_513 = {_zz_shareBuffer_sbuf_p1_rdat_514,_zz_shareBuffer_sbuf_p1_rdat_515};
  assign _zz_shareBuffer_sbuf_p1_rdat_625 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_626 = {_zz_shareBuffer_sbuf_p1_rdat_627,_zz_shareBuffer_sbuf_p1_rdat_628};
  assign _zz_shareBuffer_sbuf_p1_rdat_738 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_739 = {_zz_shareBuffer_sbuf_p1_rdat_740,_zz_shareBuffer_sbuf_p1_rdat_741};
  assign _zz_shareBuffer_sbuf_p1_rdat_851 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_852 = {_zz_shareBuffer_sbuf_p1_rdat_853,_zz_shareBuffer_sbuf_p1_rdat_854};
  assign _zz_shareBuffer_sbuf_p1_rdat_966 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_967 = {_zz_shareBuffer_sbuf_p1_rdat_968,_zz_shareBuffer_sbuf_p1_rdat_969};
  assign _zz_shareBuffer_sbuf_p1_rdat_1079 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1080 = {_zz_shareBuffer_sbuf_p1_rdat_1081,_zz_shareBuffer_sbuf_p1_rdat_1082};
  assign _zz_shareBuffer_sbuf_p1_rdat_1193 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1194 = {_zz_shareBuffer_sbuf_p1_rdat_1195,_zz_shareBuffer_sbuf_p1_rdat_1196};
  assign _zz_shareBuffer_sbuf_p1_rdat_1306 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1307 = {_zz_shareBuffer_sbuf_p1_rdat_1308,_zz_shareBuffer_sbuf_p1_rdat_1309};
  assign _zz_shareBuffer_sbuf_p1_rdat_1419 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1420 = {_zz_shareBuffer_sbuf_p1_rdat_1421,_zz_shareBuffer_sbuf_p1_rdat_1422};
  assign _zz_shareBuffer_sbuf_p1_rdat_1531 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1532 = {_zz_shareBuffer_sbuf_p1_rdat_1533,_zz_shareBuffer_sbuf_p1_rdat_1534};
  assign _zz_shareBuffer_sbuf_p1_rdat_1643 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1644 = {_zz_shareBuffer_sbuf_p1_rdat_1645,_zz_shareBuffer_sbuf_p1_rdat_1646};
  assign _zz_shareBuffer_sbuf_p1_rdat_1753 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1754 = {_zz_shareBuffer_sbuf_p1_rdat_1755,_zz_shareBuffer_sbuf_p1_rdat_1756};
  assign _zz_shareBuffer_sbuf_p1_rdat_70 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_71 = {_zz_shareBuffer_sbuf_p1_rdat_72,_zz_shareBuffer_sbuf_p1_rdat_73};
  assign _zz_shareBuffer_sbuf_p1_rdat_179 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_180 = {_zz_shareBuffer_sbuf_p1_rdat_181,_zz_shareBuffer_sbuf_p1_rdat_182};
  assign _zz_shareBuffer_sbuf_p1_rdat_290 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_291 = {_zz_shareBuffer_sbuf_p1_rdat_292,_zz_shareBuffer_sbuf_p1_rdat_293};
  assign _zz_shareBuffer_sbuf_p1_rdat_401 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_402 = {_zz_shareBuffer_sbuf_p1_rdat_403,_zz_shareBuffer_sbuf_p1_rdat_404};
  assign _zz_shareBuffer_sbuf_p1_rdat_514 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_515 = {_zz_shareBuffer_sbuf_p1_rdat_516,_zz_shareBuffer_sbuf_p1_rdat_517};
  assign _zz_shareBuffer_sbuf_p1_rdat_627 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_628 = {_zz_shareBuffer_sbuf_p1_rdat_629,_zz_shareBuffer_sbuf_p1_rdat_630};
  assign _zz_shareBuffer_sbuf_p1_rdat_740 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_741 = {_zz_shareBuffer_sbuf_p1_rdat_742,_zz_shareBuffer_sbuf_p1_rdat_743};
  assign _zz_shareBuffer_sbuf_p1_rdat_853 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_854 = {_zz_shareBuffer_sbuf_p1_rdat_855,_zz_shareBuffer_sbuf_p1_rdat_856};
  assign _zz_shareBuffer_sbuf_p1_rdat_968 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_969 = {_zz_shareBuffer_sbuf_p1_rdat_970,_zz_shareBuffer_sbuf_p1_rdat_971};
  assign _zz_shareBuffer_sbuf_p1_rdat_1081 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1082 = {_zz_shareBuffer_sbuf_p1_rdat_1083,_zz_shareBuffer_sbuf_p1_rdat_1084};
  assign _zz_shareBuffer_sbuf_p1_rdat_1195 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1196 = {_zz_shareBuffer_sbuf_p1_rdat_1197,_zz_shareBuffer_sbuf_p1_rdat_1198};
  assign _zz_shareBuffer_sbuf_p1_rdat_1308 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1309 = {_zz_shareBuffer_sbuf_p1_rdat_1310,_zz_shareBuffer_sbuf_p1_rdat_1311};
  assign _zz_shareBuffer_sbuf_p1_rdat_1421 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1422 = {_zz_shareBuffer_sbuf_p1_rdat_1423,_zz_shareBuffer_sbuf_p1_rdat_1424};
  assign _zz_shareBuffer_sbuf_p1_rdat_1533 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1534 = {_zz_shareBuffer_sbuf_p1_rdat_1535,_zz_shareBuffer_sbuf_p1_rdat_1536};
  assign _zz_shareBuffer_sbuf_p1_rdat_1645 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1646 = {_zz_shareBuffer_sbuf_p1_rdat_1647,_zz_shareBuffer_sbuf_p1_rdat_1648};
  assign _zz_shareBuffer_sbuf_p1_rdat_1755 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1756 = {_zz_shareBuffer_sbuf_p1_rdat_1757,_zz_shareBuffer_sbuf_p1_rdat_1758};
  assign _zz_shareBuffer_sbuf_p1_rdat_72 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_73 = {_zz_shareBuffer_sbuf_p1_rdat_74,_zz_shareBuffer_sbuf_p1_rdat_75};
  assign _zz_shareBuffer_sbuf_p1_rdat_181 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_182 = {_zz_shareBuffer_sbuf_p1_rdat_183,_zz_shareBuffer_sbuf_p1_rdat_184};
  assign _zz_shareBuffer_sbuf_p1_rdat_292 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_293 = {_zz_shareBuffer_sbuf_p1_rdat_294,_zz_shareBuffer_sbuf_p1_rdat_295};
  assign _zz_shareBuffer_sbuf_p1_rdat_403 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_404 = {_zz_shareBuffer_sbuf_p1_rdat_405,_zz_shareBuffer_sbuf_p1_rdat_406};
  assign _zz_shareBuffer_sbuf_p1_rdat_516 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_517 = {_zz_shareBuffer_sbuf_p1_rdat_518,_zz_shareBuffer_sbuf_p1_rdat_519};
  assign _zz_shareBuffer_sbuf_p1_rdat_629 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_630 = {_zz_shareBuffer_sbuf_p1_rdat_631,_zz_shareBuffer_sbuf_p1_rdat_632};
  assign _zz_shareBuffer_sbuf_p1_rdat_742 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_743 = {_zz_shareBuffer_sbuf_p1_rdat_744,_zz_shareBuffer_sbuf_p1_rdat_745};
  assign _zz_shareBuffer_sbuf_p1_rdat_855 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_856 = {_zz_shareBuffer_sbuf_p1_rdat_857,_zz_shareBuffer_sbuf_p1_rdat_858};
  assign _zz_shareBuffer_sbuf_p1_rdat_970 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_971 = {_zz_shareBuffer_sbuf_p1_rdat_972,_zz_shareBuffer_sbuf_p1_rdat_973};
  assign _zz_shareBuffer_sbuf_p1_rdat_1083 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1084 = {_zz_shareBuffer_sbuf_p1_rdat_1085,_zz_shareBuffer_sbuf_p1_rdat_1086};
  assign _zz_shareBuffer_sbuf_p1_rdat_1197 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1198 = {_zz_shareBuffer_sbuf_p1_rdat_1199,_zz_shareBuffer_sbuf_p1_rdat_1200};
  assign _zz_shareBuffer_sbuf_p1_rdat_1310 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1311 = {_zz_shareBuffer_sbuf_p1_rdat_1312,_zz_shareBuffer_sbuf_p1_rdat_1313};
  assign _zz_shareBuffer_sbuf_p1_rdat_1423 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1424 = {_zz_shareBuffer_sbuf_p1_rdat_1425,_zz_shareBuffer_sbuf_p1_rdat_1426};
  assign _zz_shareBuffer_sbuf_p1_rdat_1535 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1536 = {_zz_shareBuffer_sbuf_p1_rdat_1537,_zz_shareBuffer_sbuf_p1_rdat_1538};
  assign _zz_shareBuffer_sbuf_p1_rdat_1647 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1648 = {_zz_shareBuffer_sbuf_p1_rdat_1649,_zz_shareBuffer_sbuf_p1_rdat_1650};
  assign _zz_shareBuffer_sbuf_p1_rdat_1757 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1758 = {_zz_shareBuffer_sbuf_p1_rdat_1759,_zz_shareBuffer_sbuf_p1_rdat_1760};
  assign _zz_shareBuffer_sbuf_p1_rdat_74 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_75 = {_zz_shareBuffer_sbuf_p1_rdat_76,_zz_shareBuffer_sbuf_p1_rdat_77};
  assign _zz_shareBuffer_sbuf_p1_rdat_183 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_184 = {_zz_shareBuffer_sbuf_p1_rdat_185,_zz_shareBuffer_sbuf_p1_rdat_186};
  assign _zz_shareBuffer_sbuf_p1_rdat_294 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_295 = {_zz_shareBuffer_sbuf_p1_rdat_296,_zz_shareBuffer_sbuf_p1_rdat_297};
  assign _zz_shareBuffer_sbuf_p1_rdat_405 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_406 = {_zz_shareBuffer_sbuf_p1_rdat_407,_zz_shareBuffer_sbuf_p1_rdat_408};
  assign _zz_shareBuffer_sbuf_p1_rdat_518 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_519 = {_zz_shareBuffer_sbuf_p1_rdat_520,_zz_shareBuffer_sbuf_p1_rdat_521};
  assign _zz_shareBuffer_sbuf_p1_rdat_631 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_632 = {_zz_shareBuffer_sbuf_p1_rdat_633,_zz_shareBuffer_sbuf_p1_rdat_634};
  assign _zz_shareBuffer_sbuf_p1_rdat_744 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_745 = {_zz_shareBuffer_sbuf_p1_rdat_746,_zz_shareBuffer_sbuf_p1_rdat_747};
  assign _zz_shareBuffer_sbuf_p1_rdat_857 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_858 = {_zz_shareBuffer_sbuf_p1_rdat_859,_zz_shareBuffer_sbuf_p1_rdat_860};
  assign _zz_shareBuffer_sbuf_p1_rdat_972 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_973 = {_zz_shareBuffer_sbuf_p1_rdat_974,_zz_shareBuffer_sbuf_p1_rdat_975};
  assign _zz_shareBuffer_sbuf_p1_rdat_1085 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1086 = {_zz_shareBuffer_sbuf_p1_rdat_1087,_zz_shareBuffer_sbuf_p1_rdat_1088};
  assign _zz_shareBuffer_sbuf_p1_rdat_1199 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1200 = {_zz_shareBuffer_sbuf_p1_rdat_1201,_zz_shareBuffer_sbuf_p1_rdat_1202};
  assign _zz_shareBuffer_sbuf_p1_rdat_1312 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1313 = {_zz_shareBuffer_sbuf_p1_rdat_1314,_zz_shareBuffer_sbuf_p1_rdat_1315};
  assign _zz_shareBuffer_sbuf_p1_rdat_1425 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1426 = {_zz_shareBuffer_sbuf_p1_rdat_1427,_zz_shareBuffer_sbuf_p1_rdat_1428};
  assign _zz_shareBuffer_sbuf_p1_rdat_1537 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1538 = {_zz_shareBuffer_sbuf_p1_rdat_1539,_zz_shareBuffer_sbuf_p1_rdat_1540};
  assign _zz_shareBuffer_sbuf_p1_rdat_1649 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1650 = {_zz_shareBuffer_sbuf_p1_rdat_1651,_zz_shareBuffer_sbuf_p1_rdat_1652};
  assign _zz_shareBuffer_sbuf_p1_rdat_1759 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1760 = {_zz_shareBuffer_sbuf_p1_rdat_1761,_zz_shareBuffer_sbuf_p1_rdat_1762};
  assign _zz_shareBuffer_sbuf_p1_rdat_76 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_77 = {_zz_shareBuffer_sbuf_p1_rdat_78,_zz_shareBuffer_sbuf_p1_rdat_79};
  assign _zz_shareBuffer_sbuf_p1_rdat_185 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_186 = {_zz_shareBuffer_sbuf_p1_rdat_187,_zz_shareBuffer_sbuf_p1_rdat_188};
  assign _zz_shareBuffer_sbuf_p1_rdat_296 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_297 = {_zz_shareBuffer_sbuf_p1_rdat_298,_zz_shareBuffer_sbuf_p1_rdat_299};
  assign _zz_shareBuffer_sbuf_p1_rdat_407 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_408 = {_zz_shareBuffer_sbuf_p1_rdat_409,_zz_shareBuffer_sbuf_p1_rdat_410};
  assign _zz_shareBuffer_sbuf_p1_rdat_520 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_521 = {_zz_shareBuffer_sbuf_p1_rdat_522,_zz_shareBuffer_sbuf_p1_rdat_523};
  assign _zz_shareBuffer_sbuf_p1_rdat_633 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_634 = {_zz_shareBuffer_sbuf_p1_rdat_635,_zz_shareBuffer_sbuf_p1_rdat_636};
  assign _zz_shareBuffer_sbuf_p1_rdat_746 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_747 = {_zz_shareBuffer_sbuf_p1_rdat_748,_zz_shareBuffer_sbuf_p1_rdat_749};
  assign _zz_shareBuffer_sbuf_p1_rdat_859 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_860 = {_zz_shareBuffer_sbuf_p1_rdat_861,_zz_shareBuffer_sbuf_p1_rdat_862};
  assign _zz_shareBuffer_sbuf_p1_rdat_974 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_975 = {_zz_shareBuffer_sbuf_p1_rdat_976,_zz_shareBuffer_sbuf_p1_rdat_977};
  assign _zz_shareBuffer_sbuf_p1_rdat_1087 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1088 = {_zz_shareBuffer_sbuf_p1_rdat_1089,_zz_shareBuffer_sbuf_p1_rdat_1090};
  assign _zz_shareBuffer_sbuf_p1_rdat_1201 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1202 = {_zz_shareBuffer_sbuf_p1_rdat_1203,_zz_shareBuffer_sbuf_p1_rdat_1204};
  assign _zz_shareBuffer_sbuf_p1_rdat_1314 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1315 = {_zz_shareBuffer_sbuf_p1_rdat_1316,_zz_shareBuffer_sbuf_p1_rdat_1317};
  assign _zz_shareBuffer_sbuf_p1_rdat_1427 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1428 = {_zz_shareBuffer_sbuf_p1_rdat_1429,_zz_shareBuffer_sbuf_p1_rdat_1430};
  assign _zz_shareBuffer_sbuf_p1_rdat_1539 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1540 = {_zz_shareBuffer_sbuf_p1_rdat_1541,_zz_shareBuffer_sbuf_p1_rdat_1542};
  assign _zz_shareBuffer_sbuf_p1_rdat_1651 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1652 = {_zz_shareBuffer_sbuf_p1_rdat_1653,_zz_shareBuffer_sbuf_p1_rdat_1654};
  assign _zz_shareBuffer_sbuf_p1_rdat_1761 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1762 = {_zz_shareBuffer_sbuf_p1_rdat_1763,_zz_shareBuffer_sbuf_p1_rdat_1764};
  assign _zz_shareBuffer_sbuf_p1_rdat_78 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_79 = {_zz_shareBuffer_sbuf_p1_rdat_80,_zz_shareBuffer_sbuf_p1_rdat_81};
  assign _zz_shareBuffer_sbuf_p1_rdat_187 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_188 = {_zz_shareBuffer_sbuf_p1_rdat_189,_zz_shareBuffer_sbuf_p1_rdat_190};
  assign _zz_shareBuffer_sbuf_p1_rdat_298 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_299 = {_zz_shareBuffer_sbuf_p1_rdat_300,_zz_shareBuffer_sbuf_p1_rdat_301};
  assign _zz_shareBuffer_sbuf_p1_rdat_409 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_410 = {_zz_shareBuffer_sbuf_p1_rdat_411,_zz_shareBuffer_sbuf_p1_rdat_412};
  assign _zz_shareBuffer_sbuf_p1_rdat_522 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_523 = {_zz_shareBuffer_sbuf_p1_rdat_524,_zz_shareBuffer_sbuf_p1_rdat_525};
  assign _zz_shareBuffer_sbuf_p1_rdat_635 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_636 = {_zz_shareBuffer_sbuf_p1_rdat_637,_zz_shareBuffer_sbuf_p1_rdat_638};
  assign _zz_shareBuffer_sbuf_p1_rdat_748 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_749 = {_zz_shareBuffer_sbuf_p1_rdat_750,_zz_shareBuffer_sbuf_p1_rdat_751};
  assign _zz_shareBuffer_sbuf_p1_rdat_861 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_862 = {_zz_shareBuffer_sbuf_p1_rdat_863,_zz_shareBuffer_sbuf_p1_rdat_864};
  assign _zz_shareBuffer_sbuf_p1_rdat_976 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_977 = {_zz_shareBuffer_sbuf_p1_rdat_978,_zz_shareBuffer_sbuf_p1_rdat_979};
  assign _zz_shareBuffer_sbuf_p1_rdat_1089 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1090 = {_zz_shareBuffer_sbuf_p1_rdat_1091,_zz_shareBuffer_sbuf_p1_rdat_1092};
  assign _zz_shareBuffer_sbuf_p1_rdat_1203 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1204 = {_zz_shareBuffer_sbuf_p1_rdat_1205,_zz_shareBuffer_sbuf_p1_rdat_1206};
  assign _zz_shareBuffer_sbuf_p1_rdat_1316 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1317 = {_zz_shareBuffer_sbuf_p1_rdat_1318,_zz_shareBuffer_sbuf_p1_rdat_1319};
  assign _zz_shareBuffer_sbuf_p1_rdat_1429 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1430 = {_zz_shareBuffer_sbuf_p1_rdat_1431,_zz_shareBuffer_sbuf_p1_rdat_1432};
  assign _zz_shareBuffer_sbuf_p1_rdat_1541 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1542 = {_zz_shareBuffer_sbuf_p1_rdat_1543,_zz_shareBuffer_sbuf_p1_rdat_1544};
  assign _zz_shareBuffer_sbuf_p1_rdat_1653 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1654 = {_zz_shareBuffer_sbuf_p1_rdat_1655,_zz_shareBuffer_sbuf_p1_rdat_1656};
  assign _zz_shareBuffer_sbuf_p1_rdat_1763 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1764 = {_zz_shareBuffer_sbuf_p1_rdat_1765,_zz_shareBuffer_sbuf_p1_rdat_1766};
  assign _zz_shareBuffer_sbuf_p1_rdat_80 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_81 = {_zz_shareBuffer_sbuf_p1_rdat_82,_zz_shareBuffer_sbuf_p1_rdat_83};
  assign _zz_shareBuffer_sbuf_p1_rdat_189 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_190 = {_zz_shareBuffer_sbuf_p1_rdat_191,_zz_shareBuffer_sbuf_p1_rdat_192};
  assign _zz_shareBuffer_sbuf_p1_rdat_300 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_301 = {_zz_shareBuffer_sbuf_p1_rdat_302,_zz_shareBuffer_sbuf_p1_rdat_303};
  assign _zz_shareBuffer_sbuf_p1_rdat_411 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_412 = {_zz_shareBuffer_sbuf_p1_rdat_413,_zz_shareBuffer_sbuf_p1_rdat_414};
  assign _zz_shareBuffer_sbuf_p1_rdat_524 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_525 = {_zz_shareBuffer_sbuf_p1_rdat_526,_zz_shareBuffer_sbuf_p1_rdat_527};
  assign _zz_shareBuffer_sbuf_p1_rdat_637 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_638 = {_zz_shareBuffer_sbuf_p1_rdat_639,_zz_shareBuffer_sbuf_p1_rdat_640};
  assign _zz_shareBuffer_sbuf_p1_rdat_750 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_751 = {_zz_shareBuffer_sbuf_p1_rdat_752,_zz_shareBuffer_sbuf_p1_rdat_753};
  assign _zz_shareBuffer_sbuf_p1_rdat_863 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_864 = {_zz_shareBuffer_sbuf_p1_rdat_865,_zz_shareBuffer_sbuf_p1_rdat_866};
  assign _zz_shareBuffer_sbuf_p1_rdat_978 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_979 = {_zz_shareBuffer_sbuf_p1_rdat_980,_zz_shareBuffer_sbuf_p1_rdat_981};
  assign _zz_shareBuffer_sbuf_p1_rdat_1091 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1092 = {_zz_shareBuffer_sbuf_p1_rdat_1093,_zz_shareBuffer_sbuf_p1_rdat_1094};
  assign _zz_shareBuffer_sbuf_p1_rdat_1205 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1206 = {_zz_shareBuffer_sbuf_p1_rdat_1207,_zz_shareBuffer_sbuf_p1_rdat_1208};
  assign _zz_shareBuffer_sbuf_p1_rdat_1318 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1319 = {_zz_shareBuffer_sbuf_p1_rdat_1320,_zz_shareBuffer_sbuf_p1_rdat_1321};
  assign _zz_shareBuffer_sbuf_p1_rdat_1431 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1432 = {_zz_shareBuffer_sbuf_p1_rdat_1433,_zz_shareBuffer_sbuf_p1_rdat_1434};
  assign _zz_shareBuffer_sbuf_p1_rdat_1543 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1544 = {_zz_shareBuffer_sbuf_p1_rdat_1545,_zz_shareBuffer_sbuf_p1_rdat_1546};
  assign _zz_shareBuffer_sbuf_p1_rdat_1655 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1656 = {_zz_shareBuffer_sbuf_p1_rdat_1657,_zz_shareBuffer_sbuf_p1_rdat_1658};
  assign _zz_shareBuffer_sbuf_p1_rdat_1765 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1766 = {_zz_shareBuffer_sbuf_p1_rdat_1767,_zz_shareBuffer_sbuf_p1_rdat_1768};
  assign _zz_shareBuffer_sbuf_p1_rdat_82 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_83 = {_zz_shareBuffer_sbuf_p1_rdat_84,_zz_shareBuffer_sbuf_p1_rdat_85};
  assign _zz_shareBuffer_sbuf_p1_rdat_191 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_192 = {_zz_shareBuffer_sbuf_p1_rdat_193,_zz_shareBuffer_sbuf_p1_rdat_194};
  assign _zz_shareBuffer_sbuf_p1_rdat_302 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_303 = {_zz_shareBuffer_sbuf_p1_rdat_304,_zz_shareBuffer_sbuf_p1_rdat_305};
  assign _zz_shareBuffer_sbuf_p1_rdat_413 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_414 = {_zz_shareBuffer_sbuf_p1_rdat_415,_zz_shareBuffer_sbuf_p1_rdat_416};
  assign _zz_shareBuffer_sbuf_p1_rdat_526 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_527 = {_zz_shareBuffer_sbuf_p1_rdat_528,_zz_shareBuffer_sbuf_p1_rdat_529};
  assign _zz_shareBuffer_sbuf_p1_rdat_639 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_640 = {_zz_shareBuffer_sbuf_p1_rdat_641,_zz_shareBuffer_sbuf_p1_rdat_642};
  assign _zz_shareBuffer_sbuf_p1_rdat_752 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_753 = {_zz_shareBuffer_sbuf_p1_rdat_754,_zz_shareBuffer_sbuf_p1_rdat_755};
  assign _zz_shareBuffer_sbuf_p1_rdat_865 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_866 = {_zz_shareBuffer_sbuf_p1_rdat_867,_zz_shareBuffer_sbuf_p1_rdat_868};
  assign _zz_shareBuffer_sbuf_p1_rdat_980 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_981 = {_zz_shareBuffer_sbuf_p1_rdat_982,_zz_shareBuffer_sbuf_p1_rdat_983};
  assign _zz_shareBuffer_sbuf_p1_rdat_1093 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1094 = {_zz_shareBuffer_sbuf_p1_rdat_1095,_zz_shareBuffer_sbuf_p1_rdat_1096};
  assign _zz_shareBuffer_sbuf_p1_rdat_1207 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1208 = {_zz_shareBuffer_sbuf_p1_rdat_1209,_zz_shareBuffer_sbuf_p1_rdat_1210};
  assign _zz_shareBuffer_sbuf_p1_rdat_1320 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1321 = {_zz_shareBuffer_sbuf_p1_rdat_1322,_zz_shareBuffer_sbuf_p1_rdat_1323};
  assign _zz_shareBuffer_sbuf_p1_rdat_1433 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1434 = {_zz_shareBuffer_sbuf_p1_rdat_1435,_zz_shareBuffer_sbuf_p1_rdat_1436};
  assign _zz_shareBuffer_sbuf_p1_rdat_1545 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1546 = {_zz_shareBuffer_sbuf_p1_rdat_1547,_zz_shareBuffer_sbuf_p1_rdat_1548};
  assign _zz_shareBuffer_sbuf_p1_rdat_1657 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1658 = {_zz_shareBuffer_sbuf_p1_rdat_1659,_zz_shareBuffer_sbuf_p1_rdat_1660};
  assign _zz_shareBuffer_sbuf_p1_rdat_1767 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1768 = {_zz_shareBuffer_sbuf_p1_rdat_1769,_zz_shareBuffer_sbuf_p1_rdat_1770};
  assign _zz_shareBuffer_sbuf_p1_rdat_84 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_85 = {_zz_shareBuffer_sbuf_p1_rdat_86,_zz_shareBuffer_sbuf_p1_rdat_87};
  assign _zz_shareBuffer_sbuf_p1_rdat_193 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_194 = {_zz_shareBuffer_sbuf_p1_rdat_195,_zz_shareBuffer_sbuf_p1_rdat_196};
  assign _zz_shareBuffer_sbuf_p1_rdat_304 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_305 = {_zz_shareBuffer_sbuf_p1_rdat_306,_zz_shareBuffer_sbuf_p1_rdat_307};
  assign _zz_shareBuffer_sbuf_p1_rdat_415 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_416 = {_zz_shareBuffer_sbuf_p1_rdat_417,_zz_shareBuffer_sbuf_p1_rdat_418};
  assign _zz_shareBuffer_sbuf_p1_rdat_528 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_529 = {_zz_shareBuffer_sbuf_p1_rdat_530,_zz_shareBuffer_sbuf_p1_rdat_531};
  assign _zz_shareBuffer_sbuf_p1_rdat_641 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_642 = {_zz_shareBuffer_sbuf_p1_rdat_643,_zz_shareBuffer_sbuf_p1_rdat_644};
  assign _zz_shareBuffer_sbuf_p1_rdat_754 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_755 = {_zz_shareBuffer_sbuf_p1_rdat_756,_zz_shareBuffer_sbuf_p1_rdat_757};
  assign _zz_shareBuffer_sbuf_p1_rdat_867 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_868 = {_zz_shareBuffer_sbuf_p1_rdat_869,_zz_shareBuffer_sbuf_p1_rdat_870};
  assign _zz_shareBuffer_sbuf_p1_rdat_982 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_983 = {_zz_shareBuffer_sbuf_p1_rdat_984,_zz_shareBuffer_sbuf_p1_rdat_985};
  assign _zz_shareBuffer_sbuf_p1_rdat_1095 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1096 = {_zz_shareBuffer_sbuf_p1_rdat_1097,_zz_shareBuffer_sbuf_p1_rdat_1098};
  assign _zz_shareBuffer_sbuf_p1_rdat_1209 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1210 = {_zz_shareBuffer_sbuf_p1_rdat_1211,_zz_shareBuffer_sbuf_p1_rdat_1212};
  assign _zz_shareBuffer_sbuf_p1_rdat_1322 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1323 = {_zz_shareBuffer_sbuf_p1_rdat_1324,_zz_shareBuffer_sbuf_p1_rdat_1325};
  assign _zz_shareBuffer_sbuf_p1_rdat_1435 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1436 = {_zz_shareBuffer_sbuf_p1_rdat_1437,_zz_shareBuffer_sbuf_p1_rdat_1438};
  assign _zz_shareBuffer_sbuf_p1_rdat_1547 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1548 = {_zz_shareBuffer_sbuf_p1_rdat_1549,_zz_shareBuffer_sbuf_p1_rdat_1550};
  assign _zz_shareBuffer_sbuf_p1_rdat_1659 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1660 = {_zz_shareBuffer_sbuf_p1_rdat_1661,_zz_shareBuffer_sbuf_p1_rdat_1662};
  assign _zz_shareBuffer_sbuf_p1_rdat_1769 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1770 = {_zz_shareBuffer_sbuf_p1_rdat_1771,_zz_shareBuffer_sbuf_p1_rdat_1772};
  assign _zz_shareBuffer_sbuf_p1_rdat_86 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_87 = {_zz_shareBuffer_sbuf_p1_rdat_88,_zz_shareBuffer_sbuf_p1_rdat_89};
  assign _zz_shareBuffer_sbuf_p1_rdat_195 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_196 = {_zz_shareBuffer_sbuf_p1_rdat_197,_zz_shareBuffer_sbuf_p1_rdat_198};
  assign _zz_shareBuffer_sbuf_p1_rdat_306 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_307 = {_zz_shareBuffer_sbuf_p1_rdat_308,_zz_shareBuffer_sbuf_p1_rdat_309};
  assign _zz_shareBuffer_sbuf_p1_rdat_417 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_418 = {_zz_shareBuffer_sbuf_p1_rdat_419,_zz_shareBuffer_sbuf_p1_rdat_420};
  assign _zz_shareBuffer_sbuf_p1_rdat_530 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_531 = {_zz_shareBuffer_sbuf_p1_rdat_532,_zz_shareBuffer_sbuf_p1_rdat_533};
  assign _zz_shareBuffer_sbuf_p1_rdat_643 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_644 = {_zz_shareBuffer_sbuf_p1_rdat_645,_zz_shareBuffer_sbuf_p1_rdat_646};
  assign _zz_shareBuffer_sbuf_p1_rdat_756 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_757 = {_zz_shareBuffer_sbuf_p1_rdat_758,_zz_shareBuffer_sbuf_p1_rdat_759};
  assign _zz_shareBuffer_sbuf_p1_rdat_869 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_870 = {_zz_shareBuffer_sbuf_p1_rdat_871,_zz_shareBuffer_sbuf_p1_rdat_872};
  assign _zz_shareBuffer_sbuf_p1_rdat_984 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_985 = {_zz_shareBuffer_sbuf_p1_rdat_986,_zz_shareBuffer_sbuf_p1_rdat_987};
  assign _zz_shareBuffer_sbuf_p1_rdat_1097 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1098 = {_zz_shareBuffer_sbuf_p1_rdat_1099,_zz_shareBuffer_sbuf_p1_rdat_1100};
  assign _zz_shareBuffer_sbuf_p1_rdat_1211 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1212 = {_zz_shareBuffer_sbuf_p1_rdat_1213,_zz_shareBuffer_sbuf_p1_rdat_1214};
  assign _zz_shareBuffer_sbuf_p1_rdat_1324 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1325 = {_zz_shareBuffer_sbuf_p1_rdat_1326,_zz_shareBuffer_sbuf_p1_rdat_1327};
  assign _zz_shareBuffer_sbuf_p1_rdat_1437 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1438 = {_zz_shareBuffer_sbuf_p1_rdat_1439,_zz_shareBuffer_sbuf_p1_rdat_1440};
  assign _zz_shareBuffer_sbuf_p1_rdat_1549 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1550 = {_zz_shareBuffer_sbuf_p1_rdat_1551,_zz_shareBuffer_sbuf_p1_rdat_1552};
  assign _zz_shareBuffer_sbuf_p1_rdat_1661 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1662 = {_zz_shareBuffer_sbuf_p1_rdat_1663,_zz_shareBuffer_sbuf_p1_rdat_1664};
  assign _zz_shareBuffer_sbuf_p1_rdat_1771 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1772 = {_zz_shareBuffer_sbuf_p1_rdat_1773,_zz_shareBuffer_sbuf_p1_rdat_1774};
  assign _zz_shareBuffer_sbuf_p1_rdat_88 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_89 = {_zz_shareBuffer_sbuf_p1_rdat_90,_zz_shareBuffer_sbuf_p1_rdat_91};
  assign _zz_shareBuffer_sbuf_p1_rdat_197 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_198 = {_zz_shareBuffer_sbuf_p1_rdat_199,_zz_shareBuffer_sbuf_p1_rdat_200};
  assign _zz_shareBuffer_sbuf_p1_rdat_308 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_309 = {_zz_shareBuffer_sbuf_p1_rdat_310,_zz_shareBuffer_sbuf_p1_rdat_311};
  assign _zz_shareBuffer_sbuf_p1_rdat_419 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_420 = {_zz_shareBuffer_sbuf_p1_rdat_421,_zz_shareBuffer_sbuf_p1_rdat_422};
  assign _zz_shareBuffer_sbuf_p1_rdat_532 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_533 = {_zz_shareBuffer_sbuf_p1_rdat_534,_zz_shareBuffer_sbuf_p1_rdat_535};
  assign _zz_shareBuffer_sbuf_p1_rdat_645 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_646 = {_zz_shareBuffer_sbuf_p1_rdat_647,_zz_shareBuffer_sbuf_p1_rdat_648};
  assign _zz_shareBuffer_sbuf_p1_rdat_758 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_759 = {_zz_shareBuffer_sbuf_p1_rdat_760,_zz_shareBuffer_sbuf_p1_rdat_761};
  assign _zz_shareBuffer_sbuf_p1_rdat_871 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_872 = {_zz_shareBuffer_sbuf_p1_rdat_873,_zz_shareBuffer_sbuf_p1_rdat_874};
  assign _zz_shareBuffer_sbuf_p1_rdat_986 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_987 = {_zz_shareBuffer_sbuf_p1_rdat_988,_zz_shareBuffer_sbuf_p1_rdat_989};
  assign _zz_shareBuffer_sbuf_p1_rdat_1099 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1100 = {_zz_shareBuffer_sbuf_p1_rdat_1101,_zz_shareBuffer_sbuf_p1_rdat_1102};
  assign _zz_shareBuffer_sbuf_p1_rdat_1213 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1214 = {_zz_shareBuffer_sbuf_p1_rdat_1215,_zz_shareBuffer_sbuf_p1_rdat_1216};
  assign _zz_shareBuffer_sbuf_p1_rdat_1326 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1327 = {_zz_shareBuffer_sbuf_p1_rdat_1328,_zz_shareBuffer_sbuf_p1_rdat_1329};
  assign _zz_shareBuffer_sbuf_p1_rdat_1439 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1440 = {_zz_shareBuffer_sbuf_p1_rdat_1441,_zz_shareBuffer_sbuf_p1_rdat_1442};
  assign _zz_shareBuffer_sbuf_p1_rdat_1551 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1552 = {_zz_shareBuffer_sbuf_p1_rdat_1553,_zz_shareBuffer_sbuf_p1_rdat_1554};
  assign _zz_shareBuffer_sbuf_p1_rdat_1663 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1664 = {_zz_shareBuffer_sbuf_p1_rdat_1665,_zz_shareBuffer_sbuf_p1_rdat_1666};
  assign _zz_shareBuffer_sbuf_p1_rdat_1773 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1774 = {_zz_shareBuffer_sbuf_p1_rdat_1775,_zz_shareBuffer_sbuf_p1_rdat_1776};
  assign _zz_shareBuffer_sbuf_p1_rdat_90 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_91 = {_zz_shareBuffer_sbuf_p1_rdat_92,_zz_shareBuffer_sbuf_p1_rdat_93};
  assign _zz_shareBuffer_sbuf_p1_rdat_199 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_200 = {_zz_shareBuffer_sbuf_p1_rdat_201,_zz_shareBuffer_sbuf_p1_rdat_202};
  assign _zz_shareBuffer_sbuf_p1_rdat_310 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_311 = {_zz_shareBuffer_sbuf_p1_rdat_312,_zz_shareBuffer_sbuf_p1_rdat_313};
  assign _zz_shareBuffer_sbuf_p1_rdat_421 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_422 = {_zz_shareBuffer_sbuf_p1_rdat_423,_zz_shareBuffer_sbuf_p1_rdat_424};
  assign _zz_shareBuffer_sbuf_p1_rdat_534 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_535 = {_zz_shareBuffer_sbuf_p1_rdat_536,_zz_shareBuffer_sbuf_p1_rdat_537};
  assign _zz_shareBuffer_sbuf_p1_rdat_647 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_648 = {_zz_shareBuffer_sbuf_p1_rdat_649,_zz_shareBuffer_sbuf_p1_rdat_650};
  assign _zz_shareBuffer_sbuf_p1_rdat_760 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_761 = {_zz_shareBuffer_sbuf_p1_rdat_762,_zz_shareBuffer_sbuf_p1_rdat_763};
  assign _zz_shareBuffer_sbuf_p1_rdat_873 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_874 = {_zz_shareBuffer_sbuf_p1_rdat_875,_zz_shareBuffer_sbuf_p1_rdat_876};
  assign _zz_shareBuffer_sbuf_p1_rdat_988 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_989 = {_zz_shareBuffer_sbuf_p1_rdat_990,_zz_shareBuffer_sbuf_p1_rdat_991};
  assign _zz_shareBuffer_sbuf_p1_rdat_1101 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1102 = {_zz_shareBuffer_sbuf_p1_rdat_1103,_zz_shareBuffer_sbuf_p1_rdat_1104};
  assign _zz_shareBuffer_sbuf_p1_rdat_1215 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1216 = {_zz_shareBuffer_sbuf_p1_rdat_1217,_zz_shareBuffer_sbuf_p1_rdat_1218};
  assign _zz_shareBuffer_sbuf_p1_rdat_1328 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1329 = {_zz_shareBuffer_sbuf_p1_rdat_1330,_zz_shareBuffer_sbuf_p1_rdat_1331};
  assign _zz_shareBuffer_sbuf_p1_rdat_1441 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1442 = {_zz_shareBuffer_sbuf_p1_rdat_1443,_zz_shareBuffer_sbuf_p1_rdat_1444};
  assign _zz_shareBuffer_sbuf_p1_rdat_1553 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1554 = {_zz_shareBuffer_sbuf_p1_rdat_1555,_zz_shareBuffer_sbuf_p1_rdat_1556};
  assign _zz_shareBuffer_sbuf_p1_rdat_1665 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1666 = {_zz_shareBuffer_sbuf_p1_rdat_1667,_zz_shareBuffer_sbuf_p1_rdat_1668};
  assign _zz_shareBuffer_sbuf_p1_rdat_1775 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1776 = {_zz_shareBuffer_sbuf_p1_rdat_1777,_zz_shareBuffer_sbuf_p1_rdat_1778};
  assign _zz_shareBuffer_sbuf_p1_rdat_92 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_93 = {_zz_shareBuffer_sbuf_p1_rdat_94,_zz_shareBuffer_sbuf_p1_rdat_95};
  assign _zz_shareBuffer_sbuf_p1_rdat_201 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_202 = {_zz_shareBuffer_sbuf_p1_rdat_203,_zz_shareBuffer_sbuf_p1_rdat_204};
  assign _zz_shareBuffer_sbuf_p1_rdat_312 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_313 = {_zz_shareBuffer_sbuf_p1_rdat_314,_zz_shareBuffer_sbuf_p1_rdat_315};
  assign _zz_shareBuffer_sbuf_p1_rdat_423 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_424 = {_zz_shareBuffer_sbuf_p1_rdat_425,_zz_shareBuffer_sbuf_p1_rdat_426};
  assign _zz_shareBuffer_sbuf_p1_rdat_536 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_537 = {_zz_shareBuffer_sbuf_p1_rdat_538,_zz_shareBuffer_sbuf_p1_rdat_539};
  assign _zz_shareBuffer_sbuf_p1_rdat_649 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_650 = {_zz_shareBuffer_sbuf_p1_rdat_651,_zz_shareBuffer_sbuf_p1_rdat_652};
  assign _zz_shareBuffer_sbuf_p1_rdat_762 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_763 = {_zz_shareBuffer_sbuf_p1_rdat_764,_zz_shareBuffer_sbuf_p1_rdat_765};
  assign _zz_shareBuffer_sbuf_p1_rdat_875 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_876 = {_zz_shareBuffer_sbuf_p1_rdat_877,_zz_shareBuffer_sbuf_p1_rdat_878};
  assign _zz_shareBuffer_sbuf_p1_rdat_990 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_991 = {_zz_shareBuffer_sbuf_p1_rdat_992,_zz_shareBuffer_sbuf_p1_rdat_993};
  assign _zz_shareBuffer_sbuf_p1_rdat_1103 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1104 = {_zz_shareBuffer_sbuf_p1_rdat_1105,_zz_shareBuffer_sbuf_p1_rdat_1106};
  assign _zz_shareBuffer_sbuf_p1_rdat_1217 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1218 = {_zz_shareBuffer_sbuf_p1_rdat_1219,_zz_shareBuffer_sbuf_p1_rdat_1220};
  assign _zz_shareBuffer_sbuf_p1_rdat_1330 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1331 = {_zz_shareBuffer_sbuf_p1_rdat_1332,_zz_shareBuffer_sbuf_p1_rdat_1333};
  assign _zz_shareBuffer_sbuf_p1_rdat_1443 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1444 = {_zz_shareBuffer_sbuf_p1_rdat_1445,_zz_shareBuffer_sbuf_p1_rdat_1446};
  assign _zz_shareBuffer_sbuf_p1_rdat_1555 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1556 = {_zz_shareBuffer_sbuf_p1_rdat_1557,_zz_shareBuffer_sbuf_p1_rdat_1558};
  assign _zz_shareBuffer_sbuf_p1_rdat_1667 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1668 = {_zz_shareBuffer_sbuf_p1_rdat_1669,_zz_shareBuffer_sbuf_p1_rdat_1670};
  assign _zz_shareBuffer_sbuf_p1_rdat_1777 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1778 = {_zz_shareBuffer_sbuf_p1_rdat_1779,_zz_shareBuffer_sbuf_p1_rdat_1780};
  assign _zz_shareBuffer_sbuf_p1_rdat_94 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_95 = {_zz_shareBuffer_sbuf_p1_rdat_96,_zz_shareBuffer_sbuf_p1_rdat_97};
  assign _zz_shareBuffer_sbuf_p1_rdat_203 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_204 = {_zz_shareBuffer_sbuf_p1_rdat_205,_zz_shareBuffer_sbuf_p1_rdat_206};
  assign _zz_shareBuffer_sbuf_p1_rdat_314 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_315 = {_zz_shareBuffer_sbuf_p1_rdat_316,_zz_shareBuffer_sbuf_p1_rdat_317};
  assign _zz_shareBuffer_sbuf_p1_rdat_425 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_426 = {_zz_shareBuffer_sbuf_p1_rdat_427,_zz_shareBuffer_sbuf_p1_rdat_428};
  assign _zz_shareBuffer_sbuf_p1_rdat_538 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_539 = {_zz_shareBuffer_sbuf_p1_rdat_540,_zz_shareBuffer_sbuf_p1_rdat_541};
  assign _zz_shareBuffer_sbuf_p1_rdat_651 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_652 = {_zz_shareBuffer_sbuf_p1_rdat_653,_zz_shareBuffer_sbuf_p1_rdat_654};
  assign _zz_shareBuffer_sbuf_p1_rdat_764 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_765 = {_zz_shareBuffer_sbuf_p1_rdat_766,_zz_shareBuffer_sbuf_p1_rdat_767};
  assign _zz_shareBuffer_sbuf_p1_rdat_877 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_878 = {_zz_shareBuffer_sbuf_p1_rdat_879,_zz_shareBuffer_sbuf_p1_rdat_880};
  assign _zz_shareBuffer_sbuf_p1_rdat_992 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_993 = {_zz_shareBuffer_sbuf_p1_rdat_994,_zz_shareBuffer_sbuf_p1_rdat_995};
  assign _zz_shareBuffer_sbuf_p1_rdat_1105 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1106 = {_zz_shareBuffer_sbuf_p1_rdat_1107,_zz_shareBuffer_sbuf_p1_rdat_1108};
  assign _zz_shareBuffer_sbuf_p1_rdat_1219 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1220 = {_zz_shareBuffer_sbuf_p1_rdat_1221,_zz_shareBuffer_sbuf_p1_rdat_1222};
  assign _zz_shareBuffer_sbuf_p1_rdat_1332 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1333 = {_zz_shareBuffer_sbuf_p1_rdat_1334,_zz_shareBuffer_sbuf_p1_rdat_1335};
  assign _zz_shareBuffer_sbuf_p1_rdat_1445 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1446 = {_zz_shareBuffer_sbuf_p1_rdat_1447,_zz_shareBuffer_sbuf_p1_rdat_1448};
  assign _zz_shareBuffer_sbuf_p1_rdat_1557 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1558 = {_zz_shareBuffer_sbuf_p1_rdat_1559,_zz_shareBuffer_sbuf_p1_rdat_1560};
  assign _zz_shareBuffer_sbuf_p1_rdat_1669 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1670 = {_zz_shareBuffer_sbuf_p1_rdat_1671,_zz_shareBuffer_sbuf_p1_rdat_1672};
  assign _zz_shareBuffer_sbuf_p1_rdat_1779 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1780 = {_zz_shareBuffer_sbuf_p1_rdat_1781,_zz_shareBuffer_sbuf_p1_rdat_1782};
  assign _zz_shareBuffer_sbuf_p1_rdat_96 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_97 = {_zz_shareBuffer_sbuf_p1_rdat_98,_zz_shareBuffer_sbuf_p1_rdat_99};
  assign _zz_shareBuffer_sbuf_p1_rdat_205 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_206 = {_zz_shareBuffer_sbuf_p1_rdat_207,_zz_shareBuffer_sbuf_p1_rdat_208};
  assign _zz_shareBuffer_sbuf_p1_rdat_316 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_317 = {_zz_shareBuffer_sbuf_p1_rdat_318,_zz_shareBuffer_sbuf_p1_rdat_319};
  assign _zz_shareBuffer_sbuf_p1_rdat_427 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_428 = {_zz_shareBuffer_sbuf_p1_rdat_429,_zz_shareBuffer_sbuf_p1_rdat_430};
  assign _zz_shareBuffer_sbuf_p1_rdat_540 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_541 = {_zz_shareBuffer_sbuf_p1_rdat_542,_zz_shareBuffer_sbuf_p1_rdat_543};
  assign _zz_shareBuffer_sbuf_p1_rdat_653 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_654 = {_zz_shareBuffer_sbuf_p1_rdat_655,_zz_shareBuffer_sbuf_p1_rdat_656};
  assign _zz_shareBuffer_sbuf_p1_rdat_766 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_767 = {_zz_shareBuffer_sbuf_p1_rdat_768,_zz_shareBuffer_sbuf_p1_rdat_769};
  assign _zz_shareBuffer_sbuf_p1_rdat_879 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_880 = {_zz_shareBuffer_sbuf_p1_rdat_881,_zz_shareBuffer_sbuf_p1_rdat_882};
  assign _zz_shareBuffer_sbuf_p1_rdat_994 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_995 = {_zz_shareBuffer_sbuf_p1_rdat_996,_zz_shareBuffer_sbuf_p1_rdat_997};
  assign _zz_shareBuffer_sbuf_p1_rdat_1107 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1108 = {_zz_shareBuffer_sbuf_p1_rdat_1109,_zz_shareBuffer_sbuf_p1_rdat_1110};
  assign _zz_shareBuffer_sbuf_p1_rdat_1221 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1222 = {_zz_shareBuffer_sbuf_p1_rdat_1223,_zz_shareBuffer_sbuf_p1_rdat_1224};
  assign _zz_shareBuffer_sbuf_p1_rdat_1334 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1335 = {_zz_shareBuffer_sbuf_p1_rdat_1336,_zz_shareBuffer_sbuf_p1_rdat_1337};
  assign _zz_shareBuffer_sbuf_p1_rdat_1447 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1448 = {_zz_shareBuffer_sbuf_p1_rdat_1449,_zz_shareBuffer_sbuf_p1_rdat_1450};
  assign _zz_shareBuffer_sbuf_p1_rdat_1559 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1560 = {_zz_shareBuffer_sbuf_p1_rdat_1561,_zz_shareBuffer_sbuf_p1_rdat_1562};
  assign _zz_shareBuffer_sbuf_p1_rdat_1671 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1672 = {_zz_shareBuffer_sbuf_p1_rdat_1673,_zz_shareBuffer_sbuf_p1_rdat_1674};
  assign _zz_shareBuffer_sbuf_p1_rdat_1781 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1782 = {_zz_shareBuffer_sbuf_p1_rdat_1783,_zz_shareBuffer_sbuf_p1_rdat_1784};
  assign _zz_shareBuffer_sbuf_p1_rdat_98 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_99 = {_zz_shareBuffer_sbuf_p1_rdat_100,_zz_shareBuffer_sbuf_p1_rdat_101};
  assign _zz_shareBuffer_sbuf_p1_rdat_207 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_208 = {_zz_shareBuffer_sbuf_p1_rdat_209,_zz_shareBuffer_sbuf_p1_rdat_210};
  assign _zz_shareBuffer_sbuf_p1_rdat_318 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_319 = {_zz_shareBuffer_sbuf_p1_rdat_320,_zz_shareBuffer_sbuf_p1_rdat_321};
  assign _zz_shareBuffer_sbuf_p1_rdat_429 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_430 = {_zz_shareBuffer_sbuf_p1_rdat_431,_zz_shareBuffer_sbuf_p1_rdat_432};
  assign _zz_shareBuffer_sbuf_p1_rdat_542 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_543 = {_zz_shareBuffer_sbuf_p1_rdat_544,_zz_shareBuffer_sbuf_p1_rdat_545};
  assign _zz_shareBuffer_sbuf_p1_rdat_655 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_656 = {_zz_shareBuffer_sbuf_p1_rdat_657,_zz_shareBuffer_sbuf_p1_rdat_658};
  assign _zz_shareBuffer_sbuf_p1_rdat_768 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_769 = {_zz_shareBuffer_sbuf_p1_rdat_770,_zz_shareBuffer_sbuf_p1_rdat_771};
  assign _zz_shareBuffer_sbuf_p1_rdat_881 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_882 = {_zz_shareBuffer_sbuf_p1_rdat_883,_zz_shareBuffer_sbuf_p1_rdat_884};
  assign _zz_shareBuffer_sbuf_p1_rdat_996 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_997 = {_zz_shareBuffer_sbuf_p1_rdat_998,_zz_shareBuffer_sbuf_p1_rdat_999};
  assign _zz_shareBuffer_sbuf_p1_rdat_1109 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1110 = {_zz_shareBuffer_sbuf_p1_rdat_1111,_zz_shareBuffer_sbuf_p1_rdat_1112};
  assign _zz_shareBuffer_sbuf_p1_rdat_1223 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1224 = {_zz_shareBuffer_sbuf_p1_rdat_1225,_zz_shareBuffer_sbuf_p1_rdat_1226};
  assign _zz_shareBuffer_sbuf_p1_rdat_1336 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1337 = {_zz_shareBuffer_sbuf_p1_rdat_1338,_zz_shareBuffer_sbuf_p1_rdat_1339};
  assign _zz_shareBuffer_sbuf_p1_rdat_1449 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1450 = {_zz_shareBuffer_sbuf_p1_rdat_1451,_zz_shareBuffer_sbuf_p1_rdat_1452};
  assign _zz_shareBuffer_sbuf_p1_rdat_1561 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1562 = {_zz_shareBuffer_sbuf_p1_rdat_1563,_zz_shareBuffer_sbuf_p1_rdat_1564};
  assign _zz_shareBuffer_sbuf_p1_rdat_1673 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1674 = {_zz_shareBuffer_sbuf_p1_rdat_1675,_zz_shareBuffer_sbuf_p1_rdat_1676};
  assign _zz_shareBuffer_sbuf_p1_rdat_1783 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1784 = {_zz_shareBuffer_sbuf_p1_rdat_1785,_zz_shareBuffer_sbuf_p1_rdat_1786};
  assign _zz_shareBuffer_sbuf_p1_rdat_100 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_101 = {_zz_shareBuffer_sbuf_p1_rdat_102,_zz_shareBuffer_sbuf_p1_rdat_103};
  assign _zz_shareBuffer_sbuf_p1_rdat_209 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_210 = {_zz_shareBuffer_sbuf_p1_rdat_211,_zz_shareBuffer_sbuf_p1_rdat_212};
  assign _zz_shareBuffer_sbuf_p1_rdat_320 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_321 = {_zz_shareBuffer_sbuf_p1_rdat_322,_zz_shareBuffer_sbuf_p1_rdat_323};
  assign _zz_shareBuffer_sbuf_p1_rdat_431 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_432 = {_zz_shareBuffer_sbuf_p1_rdat_433,_zz_shareBuffer_sbuf_p1_rdat_434};
  assign _zz_shareBuffer_sbuf_p1_rdat_544 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_545 = {_zz_shareBuffer_sbuf_p1_rdat_546,_zz_shareBuffer_sbuf_p1_rdat_547};
  assign _zz_shareBuffer_sbuf_p1_rdat_657 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_658 = {_zz_shareBuffer_sbuf_p1_rdat_659,_zz_shareBuffer_sbuf_p1_rdat_660};
  assign _zz_shareBuffer_sbuf_p1_rdat_770 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_771 = {_zz_shareBuffer_sbuf_p1_rdat_772,_zz_shareBuffer_sbuf_p1_rdat_773};
  assign _zz_shareBuffer_sbuf_p1_rdat_883 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_884 = {_zz_shareBuffer_sbuf_p1_rdat_885,_zz_shareBuffer_sbuf_p1_rdat_886};
  assign _zz_shareBuffer_sbuf_p1_rdat_998 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_999 = {_zz_shareBuffer_sbuf_p1_rdat_1000,_zz_shareBuffer_sbuf_p1_rdat_1001};
  assign _zz_shareBuffer_sbuf_p1_rdat_1111 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1112 = {_zz_shareBuffer_sbuf_p1_rdat_1113,_zz_shareBuffer_sbuf_p1_rdat_1114};
  assign _zz_shareBuffer_sbuf_p1_rdat_1225 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1226 = {_zz_shareBuffer_sbuf_p1_rdat_1227,_zz_shareBuffer_sbuf_p1_rdat_1228};
  assign _zz_shareBuffer_sbuf_p1_rdat_1338 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1339 = {_zz_shareBuffer_sbuf_p1_rdat_1340,_zz_shareBuffer_sbuf_p1_rdat_1341};
  assign _zz_shareBuffer_sbuf_p1_rdat_1451 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1452 = {_zz_shareBuffer_sbuf_p1_rdat_1453,_zz_shareBuffer_sbuf_p1_rdat_1454};
  assign _zz_shareBuffer_sbuf_p1_rdat_1563 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1564 = {_zz_shareBuffer_sbuf_p1_rdat_1565,_zz_shareBuffer_sbuf_p1_rdat_1566};
  assign _zz_shareBuffer_sbuf_p1_rdat_1675 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1676 = {_zz_shareBuffer_sbuf_p1_rdat_1677,_zz_shareBuffer_sbuf_p1_rdat_1678};
  assign _zz_shareBuffer_sbuf_p1_rdat_1785 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1786 = {_zz_shareBuffer_sbuf_p1_rdat_1787,_zz_shareBuffer_sbuf_p1_rdat_1788};
  assign _zz_shareBuffer_sbuf_p1_rdat_102 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_103 = {shareBuffer_sbuf_p1_re_norm_d1_0,{_zz_shareBuffer_sbuf_p1_rdat_104,_zz_shareBuffer_sbuf_p1_rdat_105}};
  assign _zz_shareBuffer_sbuf_p1_rdat_211 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_212 = {shareBuffer_sbuf_p1_re_norm_d1_1,{_zz_shareBuffer_sbuf_p1_rdat_213,_zz_shareBuffer_sbuf_p1_rdat_214}};
  assign _zz_shareBuffer_sbuf_p1_rdat_322 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_323 = {shareBuffer_sbuf_p1_re_norm_d1_2,{_zz_shareBuffer_sbuf_p1_rdat_324,_zz_shareBuffer_sbuf_p1_rdat_325}};
  assign _zz_shareBuffer_sbuf_p1_rdat_433 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_434 = {shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_435,_zz_shareBuffer_sbuf_p1_rdat_436}};
  assign _zz_shareBuffer_sbuf_p1_rdat_546 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_547 = {shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_548,_zz_shareBuffer_sbuf_p1_rdat_549}};
  assign _zz_shareBuffer_sbuf_p1_rdat_659 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_660 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_661,_zz_shareBuffer_sbuf_p1_rdat_662}};
  assign _zz_shareBuffer_sbuf_p1_rdat_772 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_773 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_774,_zz_shareBuffer_sbuf_p1_rdat_775}};
  assign _zz_shareBuffer_sbuf_p1_rdat_885 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_886 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_887,_zz_shareBuffer_sbuf_p1_rdat_888}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1000 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_1001 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_1002,_zz_shareBuffer_sbuf_p1_rdat_1003}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1113 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1114 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1115,_zz_shareBuffer_sbuf_p1_rdat_1116}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1227 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1228 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1229,_zz_shareBuffer_sbuf_p1_rdat_1230}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1340 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1341 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1342,_zz_shareBuffer_sbuf_p1_rdat_1343}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1453 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1454 = {shareBuffer_sbuf_p1_re_norm_d1_12,{_zz_shareBuffer_sbuf_p1_rdat_1455,_zz_shareBuffer_sbuf_p1_rdat_1456}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1565 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1566 = {shareBuffer_sbuf_p1_re_norm_d1_13,{_zz_shareBuffer_sbuf_p1_rdat_1567,_zz_shareBuffer_sbuf_p1_rdat_1568}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1677 = shareBuffer_sbuf_p1_re_norm_d1_14;
  assign _zz_shareBuffer_sbuf_p1_rdat_1678 = {shareBuffer_sbuf_p1_re_norm_d1_14,shareBuffer_sbuf_p1_re_norm_d1_14};
  assign _zz_shareBuffer_sbuf_p1_rdat_1787 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_1788 = shareBuffer_sbuf_p1_re_norm_d1_15;
  assign _zz_shareBuffer_sbuf_p1_rdat_104 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_105 = {shareBuffer_sbuf_p1_re_norm_d1_0,{_zz_shareBuffer_sbuf_p1_rdat_106,_zz_shareBuffer_sbuf_p1_rdat_107}};
  assign _zz_shareBuffer_sbuf_p1_rdat_213 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_214 = {shareBuffer_sbuf_p1_re_norm_d1_1,{_zz_shareBuffer_sbuf_p1_rdat_215,_zz_shareBuffer_sbuf_p1_rdat_216}};
  assign _zz_shareBuffer_sbuf_p1_rdat_324 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_325 = {shareBuffer_sbuf_p1_re_norm_d1_2,{_zz_shareBuffer_sbuf_p1_rdat_326,_zz_shareBuffer_sbuf_p1_rdat_327}};
  assign _zz_shareBuffer_sbuf_p1_rdat_435 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_436 = {shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_437,_zz_shareBuffer_sbuf_p1_rdat_438}};
  assign _zz_shareBuffer_sbuf_p1_rdat_548 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_549 = {shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_550,_zz_shareBuffer_sbuf_p1_rdat_551}};
  assign _zz_shareBuffer_sbuf_p1_rdat_661 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_662 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_663,_zz_shareBuffer_sbuf_p1_rdat_664}};
  assign _zz_shareBuffer_sbuf_p1_rdat_774 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_775 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_776,_zz_shareBuffer_sbuf_p1_rdat_777}};
  assign _zz_shareBuffer_sbuf_p1_rdat_887 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_888 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_889,_zz_shareBuffer_sbuf_p1_rdat_890}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1002 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_1003 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_1004,_zz_shareBuffer_sbuf_p1_rdat_1005}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1115 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1116 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1117,_zz_shareBuffer_sbuf_p1_rdat_1118}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1229 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1230 = {shareBuffer_sbuf_p1_re_norm_d1_10,{_zz_shareBuffer_sbuf_p1_rdat_1231,_zz_shareBuffer_sbuf_p1_rdat_1232}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1342 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1343 = {shareBuffer_sbuf_p1_re_norm_d1_11,{_zz_shareBuffer_sbuf_p1_rdat_1344,_zz_shareBuffer_sbuf_p1_rdat_1345}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1455 = shareBuffer_sbuf_p1_re_norm_d1_12;
  assign _zz_shareBuffer_sbuf_p1_rdat_1456 = {shareBuffer_sbuf_p1_re_norm_d1_12,shareBuffer_sbuf_p1_re_norm_d1_12};
  assign _zz_shareBuffer_sbuf_p1_rdat_1567 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_1568 = shareBuffer_sbuf_p1_re_norm_d1_13;
  assign _zz_shareBuffer_sbuf_p1_rdat_106 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_107 = {shareBuffer_sbuf_p1_re_norm_d1_0,{_zz_shareBuffer_sbuf_p1_rdat_108,_zz_shareBuffer_sbuf_p1_rdat_109}};
  assign _zz_shareBuffer_sbuf_p1_rdat_215 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_216 = {shareBuffer_sbuf_p1_re_norm_d1_1,{_zz_shareBuffer_sbuf_p1_rdat_217,_zz_shareBuffer_sbuf_p1_rdat_218}};
  assign _zz_shareBuffer_sbuf_p1_rdat_326 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_327 = {shareBuffer_sbuf_p1_re_norm_d1_2,{_zz_shareBuffer_sbuf_p1_rdat_328,_zz_shareBuffer_sbuf_p1_rdat_329}};
  assign _zz_shareBuffer_sbuf_p1_rdat_437 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_438 = {shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_439,_zz_shareBuffer_sbuf_p1_rdat_440}};
  assign _zz_shareBuffer_sbuf_p1_rdat_550 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_551 = {shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_552,_zz_shareBuffer_sbuf_p1_rdat_553}};
  assign _zz_shareBuffer_sbuf_p1_rdat_663 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_664 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_665,_zz_shareBuffer_sbuf_p1_rdat_666}};
  assign _zz_shareBuffer_sbuf_p1_rdat_776 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_777 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_778,_zz_shareBuffer_sbuf_p1_rdat_779}};
  assign _zz_shareBuffer_sbuf_p1_rdat_889 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_890 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_891,_zz_shareBuffer_sbuf_p1_rdat_892}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1004 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_1005 = {shareBuffer_sbuf_p1_re_norm_d1_8,{_zz_shareBuffer_sbuf_p1_rdat_1006,_zz_shareBuffer_sbuf_p1_rdat_1007}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1117 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1118 = {shareBuffer_sbuf_p1_re_norm_d1_9,{_zz_shareBuffer_sbuf_p1_rdat_1119,_zz_shareBuffer_sbuf_p1_rdat_1120}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1231 = shareBuffer_sbuf_p1_re_norm_d1_10;
  assign _zz_shareBuffer_sbuf_p1_rdat_1232 = {shareBuffer_sbuf_p1_re_norm_d1_10,shareBuffer_sbuf_p1_re_norm_d1_10};
  assign _zz_shareBuffer_sbuf_p1_rdat_1344 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_1345 = shareBuffer_sbuf_p1_re_norm_d1_11;
  assign _zz_shareBuffer_sbuf_p1_rdat_108 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_109 = {shareBuffer_sbuf_p1_re_norm_d1_0,{_zz_shareBuffer_sbuf_p1_rdat_110,_zz_shareBuffer_sbuf_p1_rdat_111}};
  assign _zz_shareBuffer_sbuf_p1_rdat_217 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_218 = {shareBuffer_sbuf_p1_re_norm_d1_1,{_zz_shareBuffer_sbuf_p1_rdat_219,_zz_shareBuffer_sbuf_p1_rdat_220}};
  assign _zz_shareBuffer_sbuf_p1_rdat_328 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_329 = {shareBuffer_sbuf_p1_re_norm_d1_2,{_zz_shareBuffer_sbuf_p1_rdat_330,_zz_shareBuffer_sbuf_p1_rdat_331}};
  assign _zz_shareBuffer_sbuf_p1_rdat_439 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_440 = {shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_441,_zz_shareBuffer_sbuf_p1_rdat_442}};
  assign _zz_shareBuffer_sbuf_p1_rdat_552 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_553 = {shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_554,_zz_shareBuffer_sbuf_p1_rdat_555}};
  assign _zz_shareBuffer_sbuf_p1_rdat_665 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_666 = {shareBuffer_sbuf_p1_re_norm_d1_5,{_zz_shareBuffer_sbuf_p1_rdat_667,_zz_shareBuffer_sbuf_p1_rdat_668}};
  assign _zz_shareBuffer_sbuf_p1_rdat_778 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_779 = {shareBuffer_sbuf_p1_re_norm_d1_6,{_zz_shareBuffer_sbuf_p1_rdat_780,_zz_shareBuffer_sbuf_p1_rdat_781}};
  assign _zz_shareBuffer_sbuf_p1_rdat_891 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_892 = {shareBuffer_sbuf_p1_re_norm_d1_7,{_zz_shareBuffer_sbuf_p1_rdat_893,_zz_shareBuffer_sbuf_p1_rdat_894}};
  assign _zz_shareBuffer_sbuf_p1_rdat_1006 = shareBuffer_sbuf_p1_re_norm_d1_8;
  assign _zz_shareBuffer_sbuf_p1_rdat_1007 = {shareBuffer_sbuf_p1_re_norm_d1_8,shareBuffer_sbuf_p1_re_norm_d1_8};
  assign _zz_shareBuffer_sbuf_p1_rdat_1119 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_1120 = shareBuffer_sbuf_p1_re_norm_d1_9;
  assign _zz_shareBuffer_sbuf_p1_rdat_110 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_111 = {shareBuffer_sbuf_p1_re_norm_d1_0,{shareBuffer_sbuf_p1_re_norm_d1_0,{_zz_shareBuffer_sbuf_p1_rdat_112,_zz_shareBuffer_sbuf_p1_rdat_113}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_219 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_220 = {shareBuffer_sbuf_p1_re_norm_d1_1,{shareBuffer_sbuf_p1_re_norm_d1_1,{_zz_shareBuffer_sbuf_p1_rdat_221,_zz_shareBuffer_sbuf_p1_rdat_222}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_330 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_331 = {shareBuffer_sbuf_p1_re_norm_d1_2,{shareBuffer_sbuf_p1_re_norm_d1_2,{_zz_shareBuffer_sbuf_p1_rdat_332,_zz_shareBuffer_sbuf_p1_rdat_333}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_441 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_442 = {shareBuffer_sbuf_p1_re_norm_d1_3,{shareBuffer_sbuf_p1_re_norm_d1_3,{_zz_shareBuffer_sbuf_p1_rdat_443,_zz_shareBuffer_sbuf_p1_rdat_444}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_554 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_555 = {shareBuffer_sbuf_p1_re_norm_d1_4,{shareBuffer_sbuf_p1_re_norm_d1_4,{_zz_shareBuffer_sbuf_p1_rdat_556,_zz_shareBuffer_sbuf_p1_rdat_557}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_667 = shareBuffer_sbuf_p1_re_norm_d1_5;
  assign _zz_shareBuffer_sbuf_p1_rdat_668 = {shareBuffer_sbuf_p1_re_norm_d1_5,{shareBuffer_sbuf_p1_re_norm_d1_5,shareBuffer_sbuf_p1_re_norm_d1_5}};
  assign _zz_shareBuffer_sbuf_p1_rdat_780 = shareBuffer_sbuf_p1_re_norm_d1_6;
  assign _zz_shareBuffer_sbuf_p1_rdat_781 = {shareBuffer_sbuf_p1_re_norm_d1_6,shareBuffer_sbuf_p1_re_norm_d1_6};
  assign _zz_shareBuffer_sbuf_p1_rdat_893 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_894 = shareBuffer_sbuf_p1_re_norm_d1_7;
  assign _zz_shareBuffer_sbuf_p1_rdat_112 = shareBuffer_sbuf_p1_re_norm_d1_0;
  assign _zz_shareBuffer_sbuf_p1_rdat_113 = {shareBuffer_sbuf_p1_re_norm_d1_0,{shareBuffer_sbuf_p1_re_norm_d1_0,{shareBuffer_sbuf_p1_re_norm_d1_0,shareBuffer_sbuf_p1_re_norm_d1_0}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_221 = shareBuffer_sbuf_p1_re_norm_d1_1;
  assign _zz_shareBuffer_sbuf_p1_rdat_222 = {shareBuffer_sbuf_p1_re_norm_d1_1,{shareBuffer_sbuf_p1_re_norm_d1_1,{shareBuffer_sbuf_p1_re_norm_d1_1,shareBuffer_sbuf_p1_re_norm_d1_1}}};
  assign _zz_shareBuffer_sbuf_p1_rdat_332 = shareBuffer_sbuf_p1_re_norm_d1_2;
  assign _zz_shareBuffer_sbuf_p1_rdat_333 = {shareBuffer_sbuf_p1_re_norm_d1_2,{shareBuffer_sbuf_p1_re_norm_d1_2,shareBuffer_sbuf_p1_re_norm_d1_2}};
  assign _zz_shareBuffer_sbuf_p1_rdat_443 = shareBuffer_sbuf_p1_re_norm_d1_3;
  assign _zz_shareBuffer_sbuf_p1_rdat_444 = {shareBuffer_sbuf_p1_re_norm_d1_3,shareBuffer_sbuf_p1_re_norm_d1_3};
  assign _zz_shareBuffer_sbuf_p1_rdat_556 = shareBuffer_sbuf_p1_re_norm_d1_4;
  assign _zz_shareBuffer_sbuf_p1_rdat_557 = shareBuffer_sbuf_p1_re_norm_d1_4;
  nv_ram_rws shareBuffer_buffer_0 (
    .re    (sbuf_re_0                      ), //i
    .we    (sbuf_we_0                      ), //i
    .ra    (sbuf_ra_0[3:0]                 ), //i
    .wa    (sbuf_wa_0[3:0]                 ), //i
    .di    (sbuf_wdat_0[63:0]              ), //i
    .dout  (shareBuffer_buffer_0_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_1 (
    .re    (sbuf_re_1                      ), //i
    .we    (sbuf_we_1                      ), //i
    .ra    (sbuf_ra_1[3:0]                 ), //i
    .wa    (sbuf_wa_1[3:0]                 ), //i
    .di    (sbuf_wdat_1[63:0]              ), //i
    .dout  (shareBuffer_buffer_1_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_2 (
    .re    (sbuf_re_2                      ), //i
    .we    (sbuf_we_2                      ), //i
    .ra    (sbuf_ra_2[3:0]                 ), //i
    .wa    (sbuf_wa_2[3:0]                 ), //i
    .di    (sbuf_wdat_2[63:0]              ), //i
    .dout  (shareBuffer_buffer_2_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_3 (
    .re    (sbuf_re_3                      ), //i
    .we    (sbuf_we_3                      ), //i
    .ra    (sbuf_ra_3[3:0]                 ), //i
    .wa    (sbuf_wa_3[3:0]                 ), //i
    .di    (sbuf_wdat_3[63:0]              ), //i
    .dout  (shareBuffer_buffer_3_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_4 (
    .re    (sbuf_re_4                      ), //i
    .we    (sbuf_we_4                      ), //i
    .ra    (sbuf_ra_4[3:0]                 ), //i
    .wa    (sbuf_wa_4[3:0]                 ), //i
    .di    (sbuf_wdat_4[63:0]              ), //i
    .dout  (shareBuffer_buffer_4_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_5 (
    .re    (sbuf_re_5                      ), //i
    .we    (sbuf_we_5                      ), //i
    .ra    (sbuf_ra_5[3:0]                 ), //i
    .wa    (sbuf_wa_5[3:0]                 ), //i
    .di    (sbuf_wdat_5[63:0]              ), //i
    .dout  (shareBuffer_buffer_5_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_6 (
    .re    (sbuf_re_6                      ), //i
    .we    (sbuf_we_6                      ), //i
    .ra    (sbuf_ra_6[3:0]                 ), //i
    .wa    (sbuf_wa_6[3:0]                 ), //i
    .di    (sbuf_wdat_6[63:0]              ), //i
    .dout  (shareBuffer_buffer_6_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_7 (
    .re    (sbuf_re_7                      ), //i
    .we    (sbuf_we_7                      ), //i
    .ra    (sbuf_ra_7[3:0]                 ), //i
    .wa    (sbuf_wa_7[3:0]                 ), //i
    .di    (sbuf_wdat_7[63:0]              ), //i
    .dout  (shareBuffer_buffer_7_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_8 (
    .re    (sbuf_re_8                      ), //i
    .we    (sbuf_we_8                      ), //i
    .ra    (sbuf_ra_8[3:0]                 ), //i
    .wa    (sbuf_wa_8[3:0]                 ), //i
    .di    (sbuf_wdat_8[63:0]              ), //i
    .dout  (shareBuffer_buffer_8_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_9 (
    .re    (sbuf_re_9                      ), //i
    .we    (sbuf_we_9                      ), //i
    .ra    (sbuf_ra_9[3:0]                 ), //i
    .wa    (sbuf_wa_9[3:0]                 ), //i
    .di    (sbuf_wdat_9[63:0]              ), //i
    .dout  (shareBuffer_buffer_9_dout[63:0]), //o
    .clk   (clk                            ), //i
    .reset (reset                          )  //i
  );
  nv_ram_rws shareBuffer_buffer_10 (
    .re    (sbuf_re_10                      ), //i
    .we    (sbuf_we_10                      ), //i
    .ra    (sbuf_ra_10[3:0]                 ), //i
    .wa    (sbuf_wa_10[3:0]                 ), //i
    .di    (sbuf_wdat_10[63:0]              ), //i
    .dout  (shareBuffer_buffer_10_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  nv_ram_rws shareBuffer_buffer_11 (
    .re    (sbuf_re_11                      ), //i
    .we    (sbuf_we_11                      ), //i
    .ra    (sbuf_ra_11[3:0]                 ), //i
    .wa    (sbuf_wa_11[3:0]                 ), //i
    .di    (sbuf_wdat_11[63:0]              ), //i
    .dout  (shareBuffer_buffer_11_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  nv_ram_rws shareBuffer_buffer_12 (
    .re    (sbuf_re_12                      ), //i
    .we    (sbuf_we_12                      ), //i
    .ra    (sbuf_ra_12[3:0]                 ), //i
    .wa    (sbuf_wa_12[3:0]                 ), //i
    .di    (sbuf_wdat_12[63:0]              ), //i
    .dout  (shareBuffer_buffer_12_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  nv_ram_rws shareBuffer_buffer_13 (
    .re    (sbuf_re_13                      ), //i
    .we    (sbuf_we_13                      ), //i
    .ra    (sbuf_ra_13[3:0]                 ), //i
    .wa    (sbuf_wa_13[3:0]                 ), //i
    .di    (sbuf_wdat_13[63:0]              ), //i
    .dout  (shareBuffer_buffer_13_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  nv_ram_rws shareBuffer_buffer_14 (
    .re    (sbuf_re_14                      ), //i
    .we    (sbuf_we_14                      ), //i
    .ra    (sbuf_ra_14[3:0]                 ), //i
    .wa    (sbuf_wa_14[3:0]                 ), //i
    .di    (sbuf_wdat_14[63:0]              ), //i
    .dout  (shareBuffer_buffer_14_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  nv_ram_rws shareBuffer_buffer_15 (
    .re    (sbuf_re_15                      ), //i
    .we    (sbuf_we_15                      ), //i
    .ra    (sbuf_ra_15[3:0]                 ), //i
    .wa    (sbuf_wa_15[3:0]                 ), //i
    .di    (sbuf_wdat_15[63:0]              ), //i
    .dout  (shareBuffer_buffer_15_dout[63:0]), //o
    .clk   (clk                             ), //i
    .reset (reset                           )  //i
  );
  assign dc2sbuf_p0_wr_bsel = dc2sbuf_p_wr_0_addr_payload[7 : 4];
  assign img2sbuf_p0_wr_bsel = img2sbuf_p_wr_0_addr_payload[7 : 4];
  assign dc2sbuf_p1_wr_bsel = img2sbuf_p_wr_1_addr_payload[7 : 4];
  assign img2sbuf_p1_wr_bsel = img2sbuf_p_wr_1_addr_payload[7 : 4];
  assign dc2sbuf_p0_wr_sel_0 = ((dc2sbuf_p0_wr_bsel == 4'b0000) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_1 = ((dc2sbuf_p0_wr_bsel == 4'b0001) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_2 = ((dc2sbuf_p0_wr_bsel == 4'b0010) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_3 = ((dc2sbuf_p0_wr_bsel == 4'b0011) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_4 = ((dc2sbuf_p0_wr_bsel == 4'b0100) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_5 = ((dc2sbuf_p0_wr_bsel == 4'b0101) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_6 = ((dc2sbuf_p0_wr_bsel == 4'b0110) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_7 = ((dc2sbuf_p0_wr_bsel == 4'b0111) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_8 = ((dc2sbuf_p0_wr_bsel == 4'b1000) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_9 = ((dc2sbuf_p0_wr_bsel == 4'b1001) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_10 = ((dc2sbuf_p0_wr_bsel == 4'b1010) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_11 = ((dc2sbuf_p0_wr_bsel == 4'b1011) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_12 = ((dc2sbuf_p0_wr_bsel == 4'b1100) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_13 = ((dc2sbuf_p0_wr_bsel == 4'b1101) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_14 = ((dc2sbuf_p0_wr_bsel == 4'b1110) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p0_wr_sel_15 = ((dc2sbuf_p0_wr_bsel == 4'b1111) && dc2sbuf_p_wr_0_addr_valid);
  assign dc2sbuf_p1_wr_sel_0 = ((dc2sbuf_p1_wr_bsel == 4'b0000) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_1 = ((dc2sbuf_p1_wr_bsel == 4'b0001) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_2 = ((dc2sbuf_p1_wr_bsel == 4'b0010) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_3 = ((dc2sbuf_p1_wr_bsel == 4'b0011) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_4 = ((dc2sbuf_p1_wr_bsel == 4'b0100) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_5 = ((dc2sbuf_p1_wr_bsel == 4'b0101) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_6 = ((dc2sbuf_p1_wr_bsel == 4'b0110) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_7 = ((dc2sbuf_p1_wr_bsel == 4'b0111) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_8 = ((dc2sbuf_p1_wr_bsel == 4'b1000) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_9 = ((dc2sbuf_p1_wr_bsel == 4'b1001) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_10 = ((dc2sbuf_p1_wr_bsel == 4'b1010) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_11 = ((dc2sbuf_p1_wr_bsel == 4'b1011) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_12 = ((dc2sbuf_p1_wr_bsel == 4'b1100) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_13 = ((dc2sbuf_p1_wr_bsel == 4'b1101) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_14 = ((dc2sbuf_p1_wr_bsel == 4'b1110) && dc2sbuf_p_wr_1_addr_valid);
  assign dc2sbuf_p1_wr_sel_15 = ((dc2sbuf_p1_wr_bsel == 4'b1111) && dc2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p0_wr_sel_0 = ((img2sbuf_p0_wr_bsel == 4'b0000) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_1 = ((img2sbuf_p0_wr_bsel == 4'b0001) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_2 = ((img2sbuf_p0_wr_bsel == 4'b0010) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_3 = ((img2sbuf_p0_wr_bsel == 4'b0011) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_4 = ((img2sbuf_p0_wr_bsel == 4'b0100) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_5 = ((img2sbuf_p0_wr_bsel == 4'b0101) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_6 = ((img2sbuf_p0_wr_bsel == 4'b0110) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_7 = ((img2sbuf_p0_wr_bsel == 4'b0111) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_8 = ((img2sbuf_p0_wr_bsel == 4'b1000) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_9 = ((img2sbuf_p0_wr_bsel == 4'b1001) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_10 = ((img2sbuf_p0_wr_bsel == 4'b1010) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_11 = ((img2sbuf_p0_wr_bsel == 4'b1011) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_12 = ((img2sbuf_p0_wr_bsel == 4'b1100) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_13 = ((img2sbuf_p0_wr_bsel == 4'b1101) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_14 = ((img2sbuf_p0_wr_bsel == 4'b1110) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p0_wr_sel_15 = ((img2sbuf_p0_wr_bsel == 4'b1111) && img2sbuf_p_wr_0_addr_valid);
  assign img2sbuf_p1_wr_sel_0 = ((img2sbuf_p1_wr_bsel == 4'b0000) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_1 = ((img2sbuf_p1_wr_bsel == 4'b0001) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_2 = ((img2sbuf_p1_wr_bsel == 4'b0010) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_3 = ((img2sbuf_p1_wr_bsel == 4'b0011) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_4 = ((img2sbuf_p1_wr_bsel == 4'b0100) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_5 = ((img2sbuf_p1_wr_bsel == 4'b0101) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_6 = ((img2sbuf_p1_wr_bsel == 4'b0110) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_7 = ((img2sbuf_p1_wr_bsel == 4'b0111) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_8 = ((img2sbuf_p1_wr_bsel == 4'b1000) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_9 = ((img2sbuf_p1_wr_bsel == 4'b1001) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_10 = ((img2sbuf_p1_wr_bsel == 4'b1010) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_11 = ((img2sbuf_p1_wr_bsel == 4'b1011) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_12 = ((img2sbuf_p1_wr_bsel == 4'b1100) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_13 = ((img2sbuf_p1_wr_bsel == 4'b1101) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_14 = ((img2sbuf_p1_wr_bsel == 4'b1110) && img2sbuf_p_wr_1_addr_valid);
  assign img2sbuf_p1_wr_sel_15 = ((img2sbuf_p1_wr_bsel == 4'b1111) && img2sbuf_p_wr_1_addr_valid);
  assign sbuf_we_0 = (((dc2sbuf_p0_wr_sel_0 || dc2sbuf_p1_wr_sel_0) || img2sbuf_p0_wr_sel_0) || img2sbuf_p1_wr_sel_0);
  assign sbuf_we_1 = (((dc2sbuf_p0_wr_sel_1 || dc2sbuf_p1_wr_sel_1) || img2sbuf_p0_wr_sel_1) || img2sbuf_p1_wr_sel_1);
  assign sbuf_we_2 = (((dc2sbuf_p0_wr_sel_2 || dc2sbuf_p1_wr_sel_2) || img2sbuf_p0_wr_sel_2) || img2sbuf_p1_wr_sel_2);
  assign sbuf_we_3 = (((dc2sbuf_p0_wr_sel_3 || dc2sbuf_p1_wr_sel_3) || img2sbuf_p0_wr_sel_3) || img2sbuf_p1_wr_sel_3);
  assign sbuf_we_4 = (((dc2sbuf_p0_wr_sel_4 || dc2sbuf_p1_wr_sel_4) || img2sbuf_p0_wr_sel_4) || img2sbuf_p1_wr_sel_4);
  assign sbuf_we_5 = (((dc2sbuf_p0_wr_sel_5 || dc2sbuf_p1_wr_sel_5) || img2sbuf_p0_wr_sel_5) || img2sbuf_p1_wr_sel_5);
  assign sbuf_we_6 = (((dc2sbuf_p0_wr_sel_6 || dc2sbuf_p1_wr_sel_6) || img2sbuf_p0_wr_sel_6) || img2sbuf_p1_wr_sel_6);
  assign sbuf_we_7 = (((dc2sbuf_p0_wr_sel_7 || dc2sbuf_p1_wr_sel_7) || img2sbuf_p0_wr_sel_7) || img2sbuf_p1_wr_sel_7);
  assign sbuf_we_8 = (((dc2sbuf_p0_wr_sel_8 || dc2sbuf_p1_wr_sel_8) || img2sbuf_p0_wr_sel_8) || img2sbuf_p1_wr_sel_8);
  assign sbuf_we_9 = (((dc2sbuf_p0_wr_sel_9 || dc2sbuf_p1_wr_sel_9) || img2sbuf_p0_wr_sel_9) || img2sbuf_p1_wr_sel_9);
  assign sbuf_we_10 = (((dc2sbuf_p0_wr_sel_10 || dc2sbuf_p1_wr_sel_10) || img2sbuf_p0_wr_sel_10) || img2sbuf_p1_wr_sel_10);
  assign sbuf_we_11 = (((dc2sbuf_p0_wr_sel_11 || dc2sbuf_p1_wr_sel_11) || img2sbuf_p0_wr_sel_11) || img2sbuf_p1_wr_sel_11);
  assign sbuf_we_12 = (((dc2sbuf_p0_wr_sel_12 || dc2sbuf_p1_wr_sel_12) || img2sbuf_p0_wr_sel_12) || img2sbuf_p1_wr_sel_12);
  assign sbuf_we_13 = (((dc2sbuf_p0_wr_sel_13 || dc2sbuf_p1_wr_sel_13) || img2sbuf_p0_wr_sel_13) || img2sbuf_p1_wr_sel_13);
  assign sbuf_we_14 = (((dc2sbuf_p0_wr_sel_14 || dc2sbuf_p1_wr_sel_14) || img2sbuf_p0_wr_sel_14) || img2sbuf_p1_wr_sel_14);
  assign sbuf_we_15 = (((dc2sbuf_p0_wr_sel_15 || dc2sbuf_p1_wr_sel_15) || img2sbuf_p0_wr_sel_15) || img2sbuf_p1_wr_sel_15);
  assign sbuf_wa_0 = (((({_zz_sbuf_wa_0,_zz_sbuf_wa_0_1} & _zz_sbuf_wa_0_2) | ({_zz_sbuf_wa_0_3,_zz_sbuf_wa_0_4} & _zz_sbuf_wa_0_5)) | ({img2sbuf_p0_wr_sel_0,{_zz_sbuf_wa_0_6,_zz_sbuf_wa_0_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wa_0_8,_zz_sbuf_wa_0_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_1 = (((({_zz_sbuf_wa_1,_zz_sbuf_wa_1_1} & _zz_sbuf_wa_1_2) | ({_zz_sbuf_wa_1_3,_zz_sbuf_wa_1_4} & _zz_sbuf_wa_1_5)) | ({img2sbuf_p0_wr_sel_1,{_zz_sbuf_wa_1_6,_zz_sbuf_wa_1_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wa_1_8,_zz_sbuf_wa_1_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_2 = (((({_zz_sbuf_wa_2,_zz_sbuf_wa_2_1} & _zz_sbuf_wa_2_2) | ({_zz_sbuf_wa_2_3,_zz_sbuf_wa_2_4} & _zz_sbuf_wa_2_5)) | ({img2sbuf_p0_wr_sel_2,{_zz_sbuf_wa_2_6,_zz_sbuf_wa_2_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wa_2_8,_zz_sbuf_wa_2_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_3 = (((({_zz_sbuf_wa_3,_zz_sbuf_wa_3_1} & _zz_sbuf_wa_3_2) | ({_zz_sbuf_wa_3_3,_zz_sbuf_wa_3_4} & _zz_sbuf_wa_3_5)) | ({img2sbuf_p0_wr_sel_3,{_zz_sbuf_wa_3_6,_zz_sbuf_wa_3_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wa_3_8,_zz_sbuf_wa_3_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_4 = (((({_zz_sbuf_wa_4,_zz_sbuf_wa_4_1} & _zz_sbuf_wa_4_2) | ({_zz_sbuf_wa_4_3,_zz_sbuf_wa_4_4} & _zz_sbuf_wa_4_5)) | ({img2sbuf_p0_wr_sel_4,{_zz_sbuf_wa_4_6,_zz_sbuf_wa_4_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wa_4_8,_zz_sbuf_wa_4_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_5 = (((({_zz_sbuf_wa_5,_zz_sbuf_wa_5_1} & _zz_sbuf_wa_5_2) | ({_zz_sbuf_wa_5_3,_zz_sbuf_wa_5_4} & _zz_sbuf_wa_5_5)) | ({img2sbuf_p0_wr_sel_5,{_zz_sbuf_wa_5_6,_zz_sbuf_wa_5_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wa_5_8,_zz_sbuf_wa_5_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_6 = (((({_zz_sbuf_wa_6,_zz_sbuf_wa_6_1} & _zz_sbuf_wa_6_2) | ({_zz_sbuf_wa_6_3,_zz_sbuf_wa_6_4} & _zz_sbuf_wa_6_5)) | ({img2sbuf_p0_wr_sel_6,{_zz_sbuf_wa_6_6,_zz_sbuf_wa_6_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wa_6_8,_zz_sbuf_wa_6_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_7 = (((({_zz_sbuf_wa_7,_zz_sbuf_wa_7_1} & _zz_sbuf_wa_7_2) | ({_zz_sbuf_wa_7_3,_zz_sbuf_wa_7_4} & _zz_sbuf_wa_7_5)) | ({img2sbuf_p0_wr_sel_7,{_zz_sbuf_wa_7_6,_zz_sbuf_wa_7_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wa_7_8,_zz_sbuf_wa_7_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_8 = (((({_zz_sbuf_wa_8,_zz_sbuf_wa_8_1} & _zz_sbuf_wa_8_2) | ({_zz_sbuf_wa_8_3,_zz_sbuf_wa_8_4} & _zz_sbuf_wa_8_5)) | ({img2sbuf_p0_wr_sel_8,{_zz_sbuf_wa_8_6,_zz_sbuf_wa_8_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wa_8_8,_zz_sbuf_wa_8_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_9 = (((({_zz_sbuf_wa_9,_zz_sbuf_wa_9_1} & _zz_sbuf_wa_9_2) | ({_zz_sbuf_wa_9_3,_zz_sbuf_wa_9_4} & _zz_sbuf_wa_9_5)) | ({img2sbuf_p0_wr_sel_9,{_zz_sbuf_wa_9_6,_zz_sbuf_wa_9_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wa_9_8,_zz_sbuf_wa_9_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_10 = (((({_zz_sbuf_wa_10,_zz_sbuf_wa_10_1} & _zz_sbuf_wa_10_2) | ({_zz_sbuf_wa_10_3,_zz_sbuf_wa_10_4} & _zz_sbuf_wa_10_5)) | ({img2sbuf_p0_wr_sel_10,{_zz_sbuf_wa_10_6,_zz_sbuf_wa_10_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wa_10_8,_zz_sbuf_wa_10_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_11 = (((({_zz_sbuf_wa_11,_zz_sbuf_wa_11_1} & _zz_sbuf_wa_11_2) | ({_zz_sbuf_wa_11_3,_zz_sbuf_wa_11_4} & _zz_sbuf_wa_11_5)) | ({img2sbuf_p0_wr_sel_11,{_zz_sbuf_wa_11_6,_zz_sbuf_wa_11_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wa_11_8,_zz_sbuf_wa_11_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_12 = (((({_zz_sbuf_wa_12,_zz_sbuf_wa_12_1} & _zz_sbuf_wa_12_2) | ({_zz_sbuf_wa_12_3,_zz_sbuf_wa_12_4} & _zz_sbuf_wa_12_5)) | ({img2sbuf_p0_wr_sel_12,{_zz_sbuf_wa_12_6,_zz_sbuf_wa_12_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wa_12_8,_zz_sbuf_wa_12_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_13 = (((({_zz_sbuf_wa_13,_zz_sbuf_wa_13_1} & _zz_sbuf_wa_13_2) | ({_zz_sbuf_wa_13_3,_zz_sbuf_wa_13_4} & _zz_sbuf_wa_13_5)) | ({img2sbuf_p0_wr_sel_13,{_zz_sbuf_wa_13_6,_zz_sbuf_wa_13_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wa_13_8,_zz_sbuf_wa_13_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_14 = (((({_zz_sbuf_wa_14,_zz_sbuf_wa_14_1} & _zz_sbuf_wa_14_2) | ({_zz_sbuf_wa_14_3,_zz_sbuf_wa_14_4} & _zz_sbuf_wa_14_5)) | ({img2sbuf_p0_wr_sel_14,{_zz_sbuf_wa_14_6,_zz_sbuf_wa_14_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wa_14_8,_zz_sbuf_wa_14_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wa_15 = (((({_zz_sbuf_wa_15,_zz_sbuf_wa_15_1} & _zz_sbuf_wa_15_2) | ({_zz_sbuf_wa_15_3,_zz_sbuf_wa_15_4} & _zz_sbuf_wa_15_5)) | ({img2sbuf_p0_wr_sel_15,{_zz_sbuf_wa_15_6,_zz_sbuf_wa_15_7}} & img2sbuf_p_wr_0_addr_payload[3 : 0])) | ({img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wa_15_8,_zz_sbuf_wa_15_9}}} & img2sbuf_p_wr_1_addr_payload[3 : 0]));
  assign sbuf_wdat_0 = (((({dc2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0,_zz_sbuf_wdat_0_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_32,_zz_sbuf_wdat_0_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_0,{img2sbuf_p0_wr_sel_0,{_zz_sbuf_wdat_0_64,_zz_sbuf_wdat_0_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{img2sbuf_p1_wr_sel_0,{_zz_sbuf_wdat_0_94,_zz_sbuf_wdat_0_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_1 = (((({dc2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1,_zz_sbuf_wdat_1_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_32,_zz_sbuf_wdat_1_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_1,{img2sbuf_p0_wr_sel_1,{_zz_sbuf_wdat_1_64,_zz_sbuf_wdat_1_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{img2sbuf_p1_wr_sel_1,{_zz_sbuf_wdat_1_94,_zz_sbuf_wdat_1_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_2 = (((({dc2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2,_zz_sbuf_wdat_2_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_32,_zz_sbuf_wdat_2_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_2,{img2sbuf_p0_wr_sel_2,{_zz_sbuf_wdat_2_64,_zz_sbuf_wdat_2_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{img2sbuf_p1_wr_sel_2,{_zz_sbuf_wdat_2_94,_zz_sbuf_wdat_2_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_3 = (((({dc2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3,_zz_sbuf_wdat_3_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_32,_zz_sbuf_wdat_3_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_3,{img2sbuf_p0_wr_sel_3,{_zz_sbuf_wdat_3_64,_zz_sbuf_wdat_3_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{img2sbuf_p1_wr_sel_3,{_zz_sbuf_wdat_3_94,_zz_sbuf_wdat_3_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_4 = (((({dc2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4,_zz_sbuf_wdat_4_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_32,_zz_sbuf_wdat_4_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_4,{img2sbuf_p0_wr_sel_4,{_zz_sbuf_wdat_4_64,_zz_sbuf_wdat_4_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{img2sbuf_p1_wr_sel_4,{_zz_sbuf_wdat_4_94,_zz_sbuf_wdat_4_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_5 = (((({dc2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5,_zz_sbuf_wdat_5_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_32,_zz_sbuf_wdat_5_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_5,{img2sbuf_p0_wr_sel_5,{_zz_sbuf_wdat_5_64,_zz_sbuf_wdat_5_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{img2sbuf_p1_wr_sel_5,{_zz_sbuf_wdat_5_94,_zz_sbuf_wdat_5_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_6 = (((({dc2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6,_zz_sbuf_wdat_6_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_32,_zz_sbuf_wdat_6_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_6,{img2sbuf_p0_wr_sel_6,{_zz_sbuf_wdat_6_64,_zz_sbuf_wdat_6_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{img2sbuf_p1_wr_sel_6,{_zz_sbuf_wdat_6_94,_zz_sbuf_wdat_6_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_7 = (((({dc2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7,_zz_sbuf_wdat_7_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_32,_zz_sbuf_wdat_7_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_7,{img2sbuf_p0_wr_sel_7,{_zz_sbuf_wdat_7_64,_zz_sbuf_wdat_7_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{img2sbuf_p1_wr_sel_7,{_zz_sbuf_wdat_7_94,_zz_sbuf_wdat_7_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_8 = (((({dc2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8,_zz_sbuf_wdat_8_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_32,_zz_sbuf_wdat_8_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_8,{img2sbuf_p0_wr_sel_8,{_zz_sbuf_wdat_8_64,_zz_sbuf_wdat_8_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{img2sbuf_p1_wr_sel_8,{_zz_sbuf_wdat_8_94,_zz_sbuf_wdat_8_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_9 = (((({dc2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9,_zz_sbuf_wdat_9_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_32,_zz_sbuf_wdat_9_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_9,{img2sbuf_p0_wr_sel_9,{_zz_sbuf_wdat_9_64,_zz_sbuf_wdat_9_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{img2sbuf_p1_wr_sel_9,{_zz_sbuf_wdat_9_94,_zz_sbuf_wdat_9_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_10 = (((({dc2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10,_zz_sbuf_wdat_10_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_32,_zz_sbuf_wdat_10_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_10,{img2sbuf_p0_wr_sel_10,{_zz_sbuf_wdat_10_64,_zz_sbuf_wdat_10_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{img2sbuf_p1_wr_sel_10,{_zz_sbuf_wdat_10_94,_zz_sbuf_wdat_10_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_11 = (((({dc2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11,_zz_sbuf_wdat_11_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_32,_zz_sbuf_wdat_11_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_11,{img2sbuf_p0_wr_sel_11,{_zz_sbuf_wdat_11_64,_zz_sbuf_wdat_11_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{img2sbuf_p1_wr_sel_11,{_zz_sbuf_wdat_11_94,_zz_sbuf_wdat_11_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_12 = (((({dc2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12,_zz_sbuf_wdat_12_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_32,_zz_sbuf_wdat_12_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_12,{img2sbuf_p0_wr_sel_12,{_zz_sbuf_wdat_12_64,_zz_sbuf_wdat_12_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{img2sbuf_p1_wr_sel_12,{_zz_sbuf_wdat_12_94,_zz_sbuf_wdat_12_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_13 = (((({dc2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13,_zz_sbuf_wdat_13_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_32,_zz_sbuf_wdat_13_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_13,{img2sbuf_p0_wr_sel_13,{_zz_sbuf_wdat_13_64,_zz_sbuf_wdat_13_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{img2sbuf_p1_wr_sel_13,{_zz_sbuf_wdat_13_94,_zz_sbuf_wdat_13_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_14 = (((({dc2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14,_zz_sbuf_wdat_14_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_32,_zz_sbuf_wdat_14_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_14,{img2sbuf_p0_wr_sel_14,{_zz_sbuf_wdat_14_64,_zz_sbuf_wdat_14_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{img2sbuf_p1_wr_sel_14,{_zz_sbuf_wdat_14_94,_zz_sbuf_wdat_14_95}}}} & img2sbuf_p_wr_1_data));
  assign sbuf_wdat_15 = (((({dc2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15,_zz_sbuf_wdat_15_1}} & dc2sbuf_p_wr_0_data) | ({dc2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_32,_zz_sbuf_wdat_15_33}} & dc2sbuf_p_wr_1_data)) | ({img2sbuf_p0_wr_sel_15,{img2sbuf_p0_wr_sel_15,{_zz_sbuf_wdat_15_64,_zz_sbuf_wdat_15_65}}} & img2sbuf_p_wr_0_data)) | ({img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{img2sbuf_p1_wr_sel_15,{_zz_sbuf_wdat_15_94,_zz_sbuf_wdat_15_95}}}} & img2sbuf_p_wr_1_data));
  assign dc2sbuf_p0_rd_bsel = dc2sbuf_p_rd_0_addr_payload[7 : 4];
  assign img2sbuf_p0_rd_bsel = img2sbuf_p_rd_0_addr_payload[7 : 4];
  assign dc2sbuf_p1_rd_bsel = dc2sbuf_p_rd_1_addr_payload[7 : 4];
  assign img2sbuf_p1_rd_bsel = img2sbuf_p_rd_1_addr_payload[7 : 4];
  assign dc2sbuf_p0_rd_sel_0 = ((dc2sbuf_p0_rd_bsel == 4'b0000) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_1 = ((dc2sbuf_p0_rd_bsel == 4'b0001) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_2 = ((dc2sbuf_p0_rd_bsel == 4'b0010) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_3 = ((dc2sbuf_p0_rd_bsel == 4'b0011) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_4 = ((dc2sbuf_p0_rd_bsel == 4'b0100) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_5 = ((dc2sbuf_p0_rd_bsel == 4'b0101) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_6 = ((dc2sbuf_p0_rd_bsel == 4'b0110) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_7 = ((dc2sbuf_p0_rd_bsel == 4'b0111) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_8 = ((dc2sbuf_p0_rd_bsel == 4'b1000) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_9 = ((dc2sbuf_p0_rd_bsel == 4'b1001) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_10 = ((dc2sbuf_p0_rd_bsel == 4'b1010) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_11 = ((dc2sbuf_p0_rd_bsel == 4'b1011) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_12 = ((dc2sbuf_p0_rd_bsel == 4'b1100) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_13 = ((dc2sbuf_p0_rd_bsel == 4'b1101) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_14 = ((dc2sbuf_p0_rd_bsel == 4'b1110) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p0_rd_sel_15 = ((dc2sbuf_p0_rd_bsel == 4'b1111) && dc2sbuf_p_rd_0_addr_valid);
  assign dc2sbuf_p1_rd_sel_0 = ((dc2sbuf_p1_rd_bsel == 4'b0000) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_1 = ((dc2sbuf_p1_rd_bsel == 4'b0001) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_2 = ((dc2sbuf_p1_rd_bsel == 4'b0010) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_3 = ((dc2sbuf_p1_rd_bsel == 4'b0011) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_4 = ((dc2sbuf_p1_rd_bsel == 4'b0100) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_5 = ((dc2sbuf_p1_rd_bsel == 4'b0101) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_6 = ((dc2sbuf_p1_rd_bsel == 4'b0110) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_7 = ((dc2sbuf_p1_rd_bsel == 4'b0111) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_8 = ((dc2sbuf_p1_rd_bsel == 4'b1000) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_9 = ((dc2sbuf_p1_rd_bsel == 4'b1001) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_10 = ((dc2sbuf_p1_rd_bsel == 4'b1010) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_11 = ((dc2sbuf_p1_rd_bsel == 4'b1011) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_12 = ((dc2sbuf_p1_rd_bsel == 4'b1100) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_13 = ((dc2sbuf_p1_rd_bsel == 4'b1101) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_14 = ((dc2sbuf_p1_rd_bsel == 4'b1110) && dc2sbuf_p_rd_1_addr_valid);
  assign dc2sbuf_p1_rd_sel_15 = ((dc2sbuf_p1_rd_bsel == 4'b1111) && dc2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p0_rd_sel_0 = ((img2sbuf_p0_rd_bsel == 4'b0000) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_1 = ((img2sbuf_p0_rd_bsel == 4'b0001) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_2 = ((img2sbuf_p0_rd_bsel == 4'b0010) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_3 = ((img2sbuf_p0_rd_bsel == 4'b0011) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_4 = ((img2sbuf_p0_rd_bsel == 4'b0100) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_5 = ((img2sbuf_p0_rd_bsel == 4'b0101) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_6 = ((img2sbuf_p0_rd_bsel == 4'b0110) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_7 = ((img2sbuf_p0_rd_bsel == 4'b0111) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_8 = ((img2sbuf_p0_rd_bsel == 4'b1000) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_9 = ((img2sbuf_p0_rd_bsel == 4'b1001) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_10 = ((img2sbuf_p0_rd_bsel == 4'b1010) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_11 = ((img2sbuf_p0_rd_bsel == 4'b1011) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_12 = ((img2sbuf_p0_rd_bsel == 4'b1100) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_13 = ((img2sbuf_p0_rd_bsel == 4'b1101) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_14 = ((img2sbuf_p0_rd_bsel == 4'b1110) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p0_rd_sel_15 = ((img2sbuf_p0_rd_bsel == 4'b1111) && img2sbuf_p_rd_0_addr_valid);
  assign img2sbuf_p1_rd_sel_0 = ((img2sbuf_p1_rd_bsel == 4'b0000) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_1 = ((img2sbuf_p1_rd_bsel == 4'b0001) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_2 = ((img2sbuf_p1_rd_bsel == 4'b0010) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_3 = ((img2sbuf_p1_rd_bsel == 4'b0011) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_4 = ((img2sbuf_p1_rd_bsel == 4'b0100) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_5 = ((img2sbuf_p1_rd_bsel == 4'b0101) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_6 = ((img2sbuf_p1_rd_bsel == 4'b0110) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_7 = ((img2sbuf_p1_rd_bsel == 4'b0111) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_8 = ((img2sbuf_p1_rd_bsel == 4'b1000) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_9 = ((img2sbuf_p1_rd_bsel == 4'b1001) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_10 = ((img2sbuf_p1_rd_bsel == 4'b1010) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_11 = ((img2sbuf_p1_rd_bsel == 4'b1011) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_12 = ((img2sbuf_p1_rd_bsel == 4'b1100) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_13 = ((img2sbuf_p1_rd_bsel == 4'b1101) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_14 = ((img2sbuf_p1_rd_bsel == 4'b1110) && img2sbuf_p_rd_1_addr_valid);
  assign img2sbuf_p1_rd_sel_15 = ((img2sbuf_p1_rd_bsel == 4'b1111) && img2sbuf_p_rd_1_addr_valid);
  assign sbuf_p0_re_0 = (dc2sbuf_p0_rd_sel_0 || img2sbuf_p0_rd_sel_0);
  assign sbuf_p0_re_1 = (dc2sbuf_p0_rd_sel_1 || img2sbuf_p0_rd_sel_1);
  assign sbuf_p0_re_2 = (dc2sbuf_p0_rd_sel_2 || img2sbuf_p0_rd_sel_2);
  assign sbuf_p0_re_3 = (dc2sbuf_p0_rd_sel_3 || img2sbuf_p0_rd_sel_3);
  assign sbuf_p0_re_4 = (dc2sbuf_p0_rd_sel_4 || img2sbuf_p0_rd_sel_4);
  assign sbuf_p0_re_5 = (dc2sbuf_p0_rd_sel_5 || img2sbuf_p0_rd_sel_5);
  assign sbuf_p0_re_6 = (dc2sbuf_p0_rd_sel_6 || img2sbuf_p0_rd_sel_6);
  assign sbuf_p0_re_7 = (dc2sbuf_p0_rd_sel_7 || img2sbuf_p0_rd_sel_7);
  assign sbuf_p0_re_8 = (dc2sbuf_p0_rd_sel_8 || img2sbuf_p0_rd_sel_8);
  assign sbuf_p0_re_9 = (dc2sbuf_p0_rd_sel_9 || img2sbuf_p0_rd_sel_9);
  assign sbuf_p0_re_10 = (dc2sbuf_p0_rd_sel_10 || img2sbuf_p0_rd_sel_10);
  assign sbuf_p0_re_11 = (dc2sbuf_p0_rd_sel_11 || img2sbuf_p0_rd_sel_11);
  assign sbuf_p0_re_12 = (dc2sbuf_p0_rd_sel_12 || img2sbuf_p0_rd_sel_12);
  assign sbuf_p0_re_13 = (dc2sbuf_p0_rd_sel_13 || img2sbuf_p0_rd_sel_13);
  assign sbuf_p0_re_14 = (dc2sbuf_p0_rd_sel_14 || img2sbuf_p0_rd_sel_14);
  assign sbuf_p0_re_15 = (dc2sbuf_p0_rd_sel_15 || img2sbuf_p0_rd_sel_15);
  assign sbuf_p1_re_0 = (dc2sbuf_p1_rd_sel_0 || img2sbuf_p1_rd_sel_0);
  assign sbuf_p1_re_1 = (dc2sbuf_p1_rd_sel_1 || img2sbuf_p1_rd_sel_1);
  assign sbuf_p1_re_2 = (dc2sbuf_p1_rd_sel_2 || img2sbuf_p1_rd_sel_2);
  assign sbuf_p1_re_3 = (dc2sbuf_p1_rd_sel_3 || img2sbuf_p1_rd_sel_3);
  assign sbuf_p1_re_4 = (dc2sbuf_p1_rd_sel_4 || img2sbuf_p1_rd_sel_4);
  assign sbuf_p1_re_5 = (dc2sbuf_p1_rd_sel_5 || img2sbuf_p1_rd_sel_5);
  assign sbuf_p1_re_6 = (dc2sbuf_p1_rd_sel_6 || img2sbuf_p1_rd_sel_6);
  assign sbuf_p1_re_7 = (dc2sbuf_p1_rd_sel_7 || img2sbuf_p1_rd_sel_7);
  assign sbuf_p1_re_8 = (dc2sbuf_p1_rd_sel_8 || img2sbuf_p1_rd_sel_8);
  assign sbuf_p1_re_9 = (dc2sbuf_p1_rd_sel_9 || img2sbuf_p1_rd_sel_9);
  assign sbuf_p1_re_10 = (dc2sbuf_p1_rd_sel_10 || img2sbuf_p1_rd_sel_10);
  assign sbuf_p1_re_11 = (dc2sbuf_p1_rd_sel_11 || img2sbuf_p1_rd_sel_11);
  assign sbuf_p1_re_12 = (dc2sbuf_p1_rd_sel_12 || img2sbuf_p1_rd_sel_12);
  assign sbuf_p1_re_13 = (dc2sbuf_p1_rd_sel_13 || img2sbuf_p1_rd_sel_13);
  assign sbuf_p1_re_14 = (dc2sbuf_p1_rd_sel_14 || img2sbuf_p1_rd_sel_14);
  assign sbuf_p1_re_15 = (dc2sbuf_p1_rd_sel_15 || img2sbuf_p1_rd_sel_15);
  assign sbuf_re_0 = (sbuf_p0_re_0 || sbuf_p1_re_0);
  assign sbuf_re_1 = (sbuf_p0_re_1 || sbuf_p1_re_1);
  assign sbuf_re_2 = (sbuf_p0_re_2 || sbuf_p1_re_2);
  assign sbuf_re_3 = (sbuf_p0_re_3 || sbuf_p1_re_3);
  assign sbuf_re_4 = (sbuf_p0_re_4 || sbuf_p1_re_4);
  assign sbuf_re_5 = (sbuf_p0_re_5 || sbuf_p1_re_5);
  assign sbuf_re_6 = (sbuf_p0_re_6 || sbuf_p1_re_6);
  assign sbuf_re_7 = (sbuf_p0_re_7 || sbuf_p1_re_7);
  assign sbuf_re_8 = (sbuf_p0_re_8 || sbuf_p1_re_8);
  assign sbuf_re_9 = (sbuf_p0_re_9 || sbuf_p1_re_9);
  assign sbuf_re_10 = (sbuf_p0_re_10 || sbuf_p1_re_10);
  assign sbuf_re_11 = (sbuf_p0_re_11 || sbuf_p1_re_11);
  assign sbuf_re_12 = (sbuf_p0_re_12 || sbuf_p1_re_12);
  assign sbuf_re_13 = (sbuf_p0_re_13 || sbuf_p1_re_13);
  assign sbuf_re_14 = (sbuf_p0_re_14 || sbuf_p1_re_14);
  assign sbuf_re_15 = (sbuf_p0_re_15 || sbuf_p1_re_15);
  assign sbuf_ra_0 = (((({_zz_sbuf_ra_0,_zz_sbuf_ra_0_1} & _zz_sbuf_ra_0_2) | ({_zz_sbuf_ra_0_3,_zz_sbuf_ra_0_4} & _zz_sbuf_ra_0_5)) | ({img2sbuf_p0_rd_sel_0,{_zz_sbuf_ra_0_6,_zz_sbuf_ra_0_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_0,{img2sbuf_p1_rd_sel_0,{_zz_sbuf_ra_0_8,_zz_sbuf_ra_0_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_1 = (((({_zz_sbuf_ra_1,_zz_sbuf_ra_1_1} & _zz_sbuf_ra_1_2) | ({_zz_sbuf_ra_1_3,_zz_sbuf_ra_1_4} & _zz_sbuf_ra_1_5)) | ({img2sbuf_p0_rd_sel_1,{_zz_sbuf_ra_1_6,_zz_sbuf_ra_1_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_1,{img2sbuf_p1_rd_sel_1,{_zz_sbuf_ra_1_8,_zz_sbuf_ra_1_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_2 = (((({_zz_sbuf_ra_2,_zz_sbuf_ra_2_1} & _zz_sbuf_ra_2_2) | ({_zz_sbuf_ra_2_3,_zz_sbuf_ra_2_4} & _zz_sbuf_ra_2_5)) | ({img2sbuf_p0_rd_sel_2,{_zz_sbuf_ra_2_6,_zz_sbuf_ra_2_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_2,{img2sbuf_p1_rd_sel_2,{_zz_sbuf_ra_2_8,_zz_sbuf_ra_2_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_3 = (((({_zz_sbuf_ra_3,_zz_sbuf_ra_3_1} & _zz_sbuf_ra_3_2) | ({_zz_sbuf_ra_3_3,_zz_sbuf_ra_3_4} & _zz_sbuf_ra_3_5)) | ({img2sbuf_p0_rd_sel_3,{_zz_sbuf_ra_3_6,_zz_sbuf_ra_3_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_3,{img2sbuf_p1_rd_sel_3,{_zz_sbuf_ra_3_8,_zz_sbuf_ra_3_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_4 = (((({_zz_sbuf_ra_4,_zz_sbuf_ra_4_1} & _zz_sbuf_ra_4_2) | ({_zz_sbuf_ra_4_3,_zz_sbuf_ra_4_4} & _zz_sbuf_ra_4_5)) | ({img2sbuf_p0_rd_sel_4,{_zz_sbuf_ra_4_6,_zz_sbuf_ra_4_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_4,{img2sbuf_p1_rd_sel_4,{_zz_sbuf_ra_4_8,_zz_sbuf_ra_4_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_5 = (((({_zz_sbuf_ra_5,_zz_sbuf_ra_5_1} & _zz_sbuf_ra_5_2) | ({_zz_sbuf_ra_5_3,_zz_sbuf_ra_5_4} & _zz_sbuf_ra_5_5)) | ({img2sbuf_p0_rd_sel_5,{_zz_sbuf_ra_5_6,_zz_sbuf_ra_5_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_5,{img2sbuf_p1_rd_sel_5,{_zz_sbuf_ra_5_8,_zz_sbuf_ra_5_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_6 = (((({_zz_sbuf_ra_6,_zz_sbuf_ra_6_1} & _zz_sbuf_ra_6_2) | ({_zz_sbuf_ra_6_3,_zz_sbuf_ra_6_4} & _zz_sbuf_ra_6_5)) | ({img2sbuf_p0_rd_sel_6,{_zz_sbuf_ra_6_6,_zz_sbuf_ra_6_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_6,{img2sbuf_p1_rd_sel_6,{_zz_sbuf_ra_6_8,_zz_sbuf_ra_6_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_7 = (((({_zz_sbuf_ra_7,_zz_sbuf_ra_7_1} & _zz_sbuf_ra_7_2) | ({_zz_sbuf_ra_7_3,_zz_sbuf_ra_7_4} & _zz_sbuf_ra_7_5)) | ({img2sbuf_p0_rd_sel_7,{_zz_sbuf_ra_7_6,_zz_sbuf_ra_7_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_7,{img2sbuf_p1_rd_sel_7,{_zz_sbuf_ra_7_8,_zz_sbuf_ra_7_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_8 = (((({_zz_sbuf_ra_8,_zz_sbuf_ra_8_1} & _zz_sbuf_ra_8_2) | ({_zz_sbuf_ra_8_3,_zz_sbuf_ra_8_4} & _zz_sbuf_ra_8_5)) | ({img2sbuf_p0_rd_sel_8,{_zz_sbuf_ra_8_6,_zz_sbuf_ra_8_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_8,{img2sbuf_p1_rd_sel_8,{_zz_sbuf_ra_8_8,_zz_sbuf_ra_8_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_9 = (((({_zz_sbuf_ra_9,_zz_sbuf_ra_9_1} & _zz_sbuf_ra_9_2) | ({_zz_sbuf_ra_9_3,_zz_sbuf_ra_9_4} & _zz_sbuf_ra_9_5)) | ({img2sbuf_p0_rd_sel_9,{_zz_sbuf_ra_9_6,_zz_sbuf_ra_9_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_9,{img2sbuf_p1_rd_sel_9,{_zz_sbuf_ra_9_8,_zz_sbuf_ra_9_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_10 = (((({_zz_sbuf_ra_10,_zz_sbuf_ra_10_1} & _zz_sbuf_ra_10_2) | ({_zz_sbuf_ra_10_3,_zz_sbuf_ra_10_4} & _zz_sbuf_ra_10_5)) | ({img2sbuf_p0_rd_sel_10,{_zz_sbuf_ra_10_6,_zz_sbuf_ra_10_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_10,{img2sbuf_p1_rd_sel_10,{_zz_sbuf_ra_10_8,_zz_sbuf_ra_10_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_11 = (((({_zz_sbuf_ra_11,_zz_sbuf_ra_11_1} & _zz_sbuf_ra_11_2) | ({_zz_sbuf_ra_11_3,_zz_sbuf_ra_11_4} & _zz_sbuf_ra_11_5)) | ({img2sbuf_p0_rd_sel_11,{_zz_sbuf_ra_11_6,_zz_sbuf_ra_11_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_11,{img2sbuf_p1_rd_sel_11,{_zz_sbuf_ra_11_8,_zz_sbuf_ra_11_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_12 = (((({_zz_sbuf_ra_12,_zz_sbuf_ra_12_1} & _zz_sbuf_ra_12_2) | ({_zz_sbuf_ra_12_3,_zz_sbuf_ra_12_4} & _zz_sbuf_ra_12_5)) | ({img2sbuf_p0_rd_sel_12,{_zz_sbuf_ra_12_6,_zz_sbuf_ra_12_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_12,{img2sbuf_p1_rd_sel_12,{_zz_sbuf_ra_12_8,_zz_sbuf_ra_12_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_13 = (((({_zz_sbuf_ra_13,_zz_sbuf_ra_13_1} & _zz_sbuf_ra_13_2) | ({_zz_sbuf_ra_13_3,_zz_sbuf_ra_13_4} & _zz_sbuf_ra_13_5)) | ({img2sbuf_p0_rd_sel_13,{_zz_sbuf_ra_13_6,_zz_sbuf_ra_13_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_13,{img2sbuf_p1_rd_sel_13,{_zz_sbuf_ra_13_8,_zz_sbuf_ra_13_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_14 = (((({_zz_sbuf_ra_14,_zz_sbuf_ra_14_1} & _zz_sbuf_ra_14_2) | ({_zz_sbuf_ra_14_3,_zz_sbuf_ra_14_4} & _zz_sbuf_ra_14_5)) | ({img2sbuf_p0_rd_sel_14,{_zz_sbuf_ra_14_6,_zz_sbuf_ra_14_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_14,{img2sbuf_p1_rd_sel_14,{_zz_sbuf_ra_14_8,_zz_sbuf_ra_14_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign sbuf_ra_15 = (((({_zz_sbuf_ra_15,_zz_sbuf_ra_15_1} & _zz_sbuf_ra_15_2) | ({_zz_sbuf_ra_15_3,_zz_sbuf_ra_15_4} & _zz_sbuf_ra_15_5)) | ({img2sbuf_p0_rd_sel_15,{_zz_sbuf_ra_15_6,_zz_sbuf_ra_15_7}} & img2sbuf_p_rd_0_addr_payload[3 : 0])) | ({img2sbuf_p1_rd_sel_15,{img2sbuf_p1_rd_sel_15,{_zz_sbuf_ra_15_8,_zz_sbuf_ra_15_9}}} & img2sbuf_p_rd_1_addr_payload[3 : 0]));
  assign shareBuffer_sbuf_rdat_0 = shareBuffer_buffer_0_dout;
  assign shareBuffer_sbuf_rdat_1 = shareBuffer_buffer_1_dout;
  assign shareBuffer_sbuf_rdat_2 = shareBuffer_buffer_2_dout;
  assign shareBuffer_sbuf_rdat_3 = shareBuffer_buffer_3_dout;
  assign shareBuffer_sbuf_rdat_4 = shareBuffer_buffer_4_dout;
  assign shareBuffer_sbuf_rdat_5 = shareBuffer_buffer_5_dout;
  assign shareBuffer_sbuf_rdat_6 = shareBuffer_buffer_6_dout;
  assign shareBuffer_sbuf_rdat_7 = shareBuffer_buffer_7_dout;
  assign shareBuffer_sbuf_rdat_8 = shareBuffer_buffer_8_dout;
  assign shareBuffer_sbuf_rdat_9 = shareBuffer_buffer_9_dout;
  assign shareBuffer_sbuf_rdat_10 = shareBuffer_buffer_10_dout;
  assign shareBuffer_sbuf_rdat_11 = shareBuffer_buffer_11_dout;
  assign shareBuffer_sbuf_rdat_12 = shareBuffer_buffer_12_dout;
  assign shareBuffer_sbuf_rdat_13 = shareBuffer_buffer_13_dout;
  assign shareBuffer_sbuf_rdat_14 = shareBuffer_buffer_14_dout;
  assign shareBuffer_sbuf_rdat_15 = shareBuffer_buffer_15_dout;
  assign shareBuffer_sbuf_p0_rdat = (((((_zz_shareBuffer_sbuf_p0_rdat | _zz_shareBuffer_sbuf_p0_rdat_1233) | (_zz_shareBuffer_sbuf_p0_rdat_1346 & shareBuffer_sbuf_rdat_12)) | ({_zz_shareBuffer_sbuf_p0_rdat_1457,_zz_shareBuffer_sbuf_p0_rdat_1458} & shareBuffer_sbuf_rdat_13)) | ({shareBuffer_sbuf_p0_re_norm_d1_14,{_zz_shareBuffer_sbuf_p0_rdat_1569,_zz_shareBuffer_sbuf_p0_rdat_1570}} & shareBuffer_sbuf_rdat_14)) | ({shareBuffer_sbuf_p0_re_norm_d1_15,{shareBuffer_sbuf_p0_re_norm_d1_15,{_zz_shareBuffer_sbuf_p0_rdat_1679,_zz_shareBuffer_sbuf_p0_rdat_1680}}} & shareBuffer_sbuf_rdat_15));
  assign shareBuffer_sbuf_p1_rdat = (((((_zz_shareBuffer_sbuf_p1_rdat | _zz_shareBuffer_sbuf_p1_rdat_1233) | (_zz_shareBuffer_sbuf_p1_rdat_1346 & shareBuffer_sbuf_rdat_12)) | ({_zz_shareBuffer_sbuf_p1_rdat_1457,_zz_shareBuffer_sbuf_p1_rdat_1458} & shareBuffer_sbuf_rdat_13)) | ({shareBuffer_sbuf_p1_re_norm_d1_14,{_zz_shareBuffer_sbuf_p1_rdat_1569,_zz_shareBuffer_sbuf_p1_rdat_1570}} & shareBuffer_sbuf_rdat_14)) | ({shareBuffer_sbuf_p1_re_norm_d1_15,{shareBuffer_sbuf_p1_re_norm_d1_15,{_zz_shareBuffer_sbuf_p1_rdat_1679,_zz_shareBuffer_sbuf_p1_rdat_1680}}} & shareBuffer_sbuf_rdat_15));
  assign dc2sbuf_p_rd_0_data = shareBuffer_sbuf_p0_rdat_d2;
  assign img2sbuf_p_rd_0_data = shareBuffer_sbuf_p0_rdat_d2;
  assign dc2sbuf_p_rd_1_data = shareBuffer_sbuf_p1_rdat_d2;
  assign img2sbuf_p_rd_1_data = shareBuffer_sbuf_p1_rdat_d2;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      shareBuffer_sbuf_p0_re_norm_d1_0 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_1 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_2 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_3 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_4 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_5 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_6 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_7 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_8 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_9 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_10 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_11 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_12 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_13 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_14 <= 1'b0;
      shareBuffer_sbuf_p0_re_norm_d1_15 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_0 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_1 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_2 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_3 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_4 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_5 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_6 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_7 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_8 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_9 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_10 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_11 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_12 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_13 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_14 <= 1'b0;
      shareBuffer_sbuf_p1_re_norm_d1_15 <= 1'b0;
      shareBuffer_sbuf_p0_rd_en_d1 <= 1'b0;
      shareBuffer_sbuf_p1_rd_en_d1 <= 1'b0;
    end else begin
      shareBuffer_sbuf_p0_re_norm_d1_0 <= sbuf_p0_re_0;
      shareBuffer_sbuf_p1_re_norm_d1_0 <= sbuf_p1_re_0;
      shareBuffer_sbuf_p0_re_norm_d1_1 <= sbuf_p0_re_1;
      shareBuffer_sbuf_p1_re_norm_d1_1 <= sbuf_p1_re_1;
      shareBuffer_sbuf_p0_re_norm_d1_2 <= sbuf_p0_re_2;
      shareBuffer_sbuf_p1_re_norm_d1_2 <= sbuf_p1_re_2;
      shareBuffer_sbuf_p0_re_norm_d1_3 <= sbuf_p0_re_3;
      shareBuffer_sbuf_p1_re_norm_d1_3 <= sbuf_p1_re_3;
      shareBuffer_sbuf_p0_re_norm_d1_4 <= sbuf_p0_re_4;
      shareBuffer_sbuf_p1_re_norm_d1_4 <= sbuf_p1_re_4;
      shareBuffer_sbuf_p0_re_norm_d1_5 <= sbuf_p0_re_5;
      shareBuffer_sbuf_p1_re_norm_d1_5 <= sbuf_p1_re_5;
      shareBuffer_sbuf_p0_re_norm_d1_6 <= sbuf_p0_re_6;
      shareBuffer_sbuf_p1_re_norm_d1_6 <= sbuf_p1_re_6;
      shareBuffer_sbuf_p0_re_norm_d1_7 <= sbuf_p0_re_7;
      shareBuffer_sbuf_p1_re_norm_d1_7 <= sbuf_p1_re_7;
      shareBuffer_sbuf_p0_re_norm_d1_8 <= sbuf_p0_re_8;
      shareBuffer_sbuf_p1_re_norm_d1_8 <= sbuf_p1_re_8;
      shareBuffer_sbuf_p0_re_norm_d1_9 <= sbuf_p0_re_9;
      shareBuffer_sbuf_p1_re_norm_d1_9 <= sbuf_p1_re_9;
      shareBuffer_sbuf_p0_re_norm_d1_10 <= sbuf_p0_re_10;
      shareBuffer_sbuf_p1_re_norm_d1_10 <= sbuf_p1_re_10;
      shareBuffer_sbuf_p0_re_norm_d1_11 <= sbuf_p0_re_11;
      shareBuffer_sbuf_p1_re_norm_d1_11 <= sbuf_p1_re_11;
      shareBuffer_sbuf_p0_re_norm_d1_12 <= sbuf_p0_re_12;
      shareBuffer_sbuf_p1_re_norm_d1_12 <= sbuf_p1_re_12;
      shareBuffer_sbuf_p0_re_norm_d1_13 <= sbuf_p0_re_13;
      shareBuffer_sbuf_p1_re_norm_d1_13 <= sbuf_p1_re_13;
      shareBuffer_sbuf_p0_re_norm_d1_14 <= sbuf_p0_re_14;
      shareBuffer_sbuf_p1_re_norm_d1_14 <= sbuf_p1_re_14;
      shareBuffer_sbuf_p0_re_norm_d1_15 <= sbuf_p0_re_15;
      shareBuffer_sbuf_p1_re_norm_d1_15 <= sbuf_p1_re_15;
      shareBuffer_sbuf_p0_rd_en_d1 <= (dc2sbuf_p_rd_0_addr_valid || img2sbuf_p_rd_0_addr_valid);
      shareBuffer_sbuf_p1_rd_en_d1 <= (dc2sbuf_p_rd_1_addr_valid || img2sbuf_p_rd_1_addr_valid);
    end
  end

  always @(posedge clk) begin
    if(shareBuffer_sbuf_p0_rd_en_d1) begin
      shareBuffer_sbuf_p0_rdat_d2 <= shareBuffer_sbuf_p0_rdat;
    end
    if(shareBuffer_sbuf_p1_rd_en_d1) begin
      shareBuffer_sbuf_p1_rdat_d2 <= shareBuffer_sbuf_p1_rdat;
    end
  end


endmodule

//nv_ram_rws_15 replaced by nv_ram_rws

//nv_ram_rws_14 replaced by nv_ram_rws

//nv_ram_rws_13 replaced by nv_ram_rws

//nv_ram_rws_12 replaced by nv_ram_rws

//nv_ram_rws_11 replaced by nv_ram_rws

//nv_ram_rws_10 replaced by nv_ram_rws

//nv_ram_rws_9 replaced by nv_ram_rws

//nv_ram_rws_8 replaced by nv_ram_rws

//nv_ram_rws_7 replaced by nv_ram_rws

//nv_ram_rws_6 replaced by nv_ram_rws

//nv_ram_rws_5 replaced by nv_ram_rws

//nv_ram_rws_4 replaced by nv_ram_rws

//nv_ram_rws_3 replaced by nv_ram_rws

//nv_ram_rws_2 replaced by nv_ram_rws

//nv_ram_rws_1 replaced by nv_ram_rws

module nv_ram_rws (
  input  wire          re,
  input  wire          we,
  input  wire [3:0]    ra,
  input  wire [3:0]    wa,
  input  wire [63:0]   di,
  output wire [63:0]   dout,
  input  wire          clk,
  input  wire          reset
);

  reg        [63:0]   _zz__zz_1_port1;
  reg [63:0] _zz_1 [0:15];

  always @(posedge clk) begin
    if(we) begin
      _zz_1[wa] <= di;
    end
  end

  always @(posedge clk) begin
    if(re) begin
      _zz__zz_1_port1 <= _zz_1[ra];
    end
  end

  assign dout = _zz__zz_1_port1;

endmodule
